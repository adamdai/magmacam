module main (input  CLKIN);
endmodule

