//Module: Add16 defined externally
//Module: pullresistor defined externally


module coreir_mux #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  input sel,
  output [width-1:0] out
);
  assign out = sel ? in1 : in0;

endmodule //coreir_mux

module bitopn_U19 (
  input [0:0] in,
  output  out
);
  //All the connections
  assign out = in[0];

endmodule //bitopn_U19

module coreir_const #(parameter value=1, parameter width=1) (
  output [width-1:0] out
);
  assign out = value;

endmodule //coreir_const

module corebit_and (
  input in0,
  input in1,
  output out
);
  assign out = in0 & in1;

endmodule //corebit_and

module bitopn_U18 (
  input [1:0] in,
  output  out
);
  //Wire declarations for instance 'join' (Module corebit_and)
  wire  join__in0;
  wire  join__in1;
  wire  join__out;
  corebit_and join(
    .in0(join__in0),
    .in1(join__in1),
    .out(join__out)
  );

  //All the connections
  assign join__in0 = in[0];
  assign out = join__out;
  assign join__in1 = in[1];

endmodule //bitopn_U18

module bitopn_U9 (
  input [2:0] in,
  output  out
);
  //Wire declarations for instance 'join' (Module corebit_and)
  wire  join__in0;
  wire  join__in1;
  wire  join__out;
  corebit_and join(
    .in0(join__in0),
    .in1(join__in1),
    .out(join__out)
  );

  //Wire declarations for instance 'opN_0' (Module bitopn_U18)
  wire [1:0] opN_0__in;
  wire  opN_0__out;
  bitopn_U18 opN_0(
    .in(opN_0__in),
    .out(opN_0__out)
  );

  //Wire declarations for instance 'opN_1' (Module bitopn_U19)
  wire [0:0] opN_1__in;
  wire  opN_1__out;
  bitopn_U19 opN_1(
    .in(opN_1__in),
    .out(opN_1__out)
  );

  //All the connections
  assign out = join__out;
  assign join__in0 = opN_0__out;
  assign opN_0__in[1] = in[1];
  assign opN_0__in[0] = in[0];
  assign join__in1 = opN_1__out;
  assign opN_1__in[0] = in[2];

endmodule //bitopn_U9

module corebit_concat (
  input in0,
  input in1,
  output [1:0] out
);
  assign out = {in0, in1};

endmodule //corebit_concat

module corebit_const #(parameter value=1) (
  output out
);
  assign out = value;

endmodule //corebit_const

module corebit_ibuf (
  inout in,
  output out
);
  assign out = in;

endmodule //corebit_ibuf

module corebit_mux (
  input in0,
  input in1,
  input sel,
  output out
);
  assign out = sel ? in1 : in0;

endmodule //corebit_mux

module corebit_not (
  input in,
  output out
);
  assign out = ~in;

endmodule //corebit_not

module corebit_or (
  input in0,
  input in1,
  output out
);
  assign out = in0 | in1;

endmodule //corebit_or

module corebit_reg #(parameter clk_posedge=1, parameter init=1) (
  input clk,
  input in,
  output out
);
reg outReg = init;
always @(posedge clk) begin
  outReg <= in;
end
assign out = outReg;

endmodule //corebit_reg

module coreir_add #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output [width-1:0] out
);
  assign out = in0 + in1;

endmodule //coreir_add

module corebit_reg_arst #(parameter arst_posedge=1, parameter clk_posedge=1, parameter init=1) (
  input clk,
  input in,
  input arst,
  output out
);
reg outReg;
wire real_rst;
assign real_rst = arst_posedge ? arst : ~arst;
wire real_clk;
assign real_clk = clk_posedge ? clk : ~clk;
always @(posedge real_clk, posedge real_rst) begin
  if (real_rst) outReg <= init;
  else outReg <= in;
end
assign out = outReg;

endmodule //corebit_reg_arst

module corebit_term (
  input in
);


endmodule //corebit_term

module corebit_tribuf (
  input in,
  input en,
  inout out
);
  assign out = en ? in : 1'bz;

endmodule //corebit_tribuf

module corebit_wire (
  input in,
  output out
);
  assign out = in;

endmodule //corebit_wire

module corebit_xor (
  input in0,
  input in1,
  output out
);
  assign out = in0 ^ in1;

endmodule //corebit_xor

module coreir_zext #(parameter width_in=1, parameter width_out=1) (
  input [width_in-1:0] in,
  output [width_out-1:0] out
);
  assign out = {{(width_out-width_in){1'b0}},in};

endmodule //coreir_zext

module coreir_eq #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output out
);
  assign out = in0 == in1;

endmodule //coreir_eq

module coreir_mem #(parameter depth=1, parameter has_init=1, parameter width=1) (
  input clk,
  input [width-1:0] wdata,
  input [$clog2(depth)-1:0] waddr,
  input wen,
  output [width-1:0] rdata,
  input [$clog2(depth)-1:0] raddr
);
reg [width-1:0] data[depth-1:0];
always @(posedge clk) begin
  if (wen) begin
    data[waddr] <= wdata;
  end
end
assign rdata = data[raddr];

endmodule //coreir_mem

module coreir_or #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output [width-1:0] out
);
  assign out = in0 | in1;

endmodule //coreir_or

module coreir_reg #(parameter clk_posedge=1, parameter init=1, parameter width=1) (
  input clk,
  input [width-1:0] in,
  output [width-1:0] out
);
reg [width-1:0] outReg=init;
wire real_clk;
assign real_clk = clk_posedge ? clk : ~clk;
always @(posedge real_clk) begin
  outReg <= in;
end
assign out = outReg;

endmodule //coreir_reg

module linebuffer_U3 (
  input  clk,
  input [15:0] in_0,
  output [15:0] out_0,
  output [15:0] out_1,
  output [15:0] out_10,
  output [15:0] out_11,
  output [15:0] out_12,
  output [15:0] out_13,
  output [15:0] out_14,
  output [15:0] out_15,
  output [15:0] out_16,
  output [15:0] out_17,
  output [15:0] out_18,
  output [15:0] out_19,
  output [15:0] out_2,
  output [15:0] out_3,
  output [15:0] out_4,
  output [15:0] out_5,
  output [15:0] out_6,
  output [15:0] out_7,
  output [15:0] out_8,
  output [15:0] out_9,
  output  valid,
  output  valid_chain,
  input  wen
);
  //Wire declarations for instance 'reg_1' (Module coreir_reg)
  wire  reg_1__clk;
  wire [15:0] reg_1__in;
  wire [15:0] reg_1__out;
  coreir_reg #(.clk_posedge(1),.init(16'bxxxxxxxxxxxxxxxx),.width(16)) reg_1(
    .clk(reg_1__clk),
    .in(reg_1__in),
    .out(reg_1__out)
  );

  //Wire declarations for instance 'reg_10' (Module coreir_reg)
  wire  reg_10__clk;
  wire [15:0] reg_10__in;
  wire [15:0] reg_10__out;
  coreir_reg #(.clk_posedge(1),.init(16'bxxxxxxxxxxxxxxxx),.width(16)) reg_10(
    .clk(reg_10__clk),
    .in(reg_10__in),
    .out(reg_10__out)
  );

  //Wire declarations for instance 'reg_11' (Module coreir_reg)
  wire  reg_11__clk;
  wire [15:0] reg_11__in;
  wire [15:0] reg_11__out;
  coreir_reg #(.clk_posedge(1),.init(16'bxxxxxxxxxxxxxxxx),.width(16)) reg_11(
    .clk(reg_11__clk),
    .in(reg_11__in),
    .out(reg_11__out)
  );

  //Wire declarations for instance 'reg_12' (Module coreir_reg)
  wire  reg_12__clk;
  wire [15:0] reg_12__in;
  wire [15:0] reg_12__out;
  coreir_reg #(.clk_posedge(1),.init(16'bxxxxxxxxxxxxxxxx),.width(16)) reg_12(
    .clk(reg_12__clk),
    .in(reg_12__in),
    .out(reg_12__out)
  );

  //Wire declarations for instance 'reg_13' (Module coreir_reg)
  wire  reg_13__clk;
  wire [15:0] reg_13__in;
  wire [15:0] reg_13__out;
  coreir_reg #(.clk_posedge(1),.init(16'bxxxxxxxxxxxxxxxx),.width(16)) reg_13(
    .clk(reg_13__clk),
    .in(reg_13__in),
    .out(reg_13__out)
  );

  //Wire declarations for instance 'reg_14' (Module coreir_reg)
  wire  reg_14__clk;
  wire [15:0] reg_14__in;
  wire [15:0] reg_14__out;
  coreir_reg #(.clk_posedge(1),.init(16'bxxxxxxxxxxxxxxxx),.width(16)) reg_14(
    .clk(reg_14__clk),
    .in(reg_14__in),
    .out(reg_14__out)
  );

  //Wire declarations for instance 'reg_15' (Module coreir_reg)
  wire  reg_15__clk;
  wire [15:0] reg_15__in;
  wire [15:0] reg_15__out;
  coreir_reg #(.clk_posedge(1),.init(16'bxxxxxxxxxxxxxxxx),.width(16)) reg_15(
    .clk(reg_15__clk),
    .in(reg_15__in),
    .out(reg_15__out)
  );

  //Wire declarations for instance 'reg_16' (Module coreir_reg)
  wire  reg_16__clk;
  wire [15:0] reg_16__in;
  wire [15:0] reg_16__out;
  coreir_reg #(.clk_posedge(1),.init(16'bxxxxxxxxxxxxxxxx),.width(16)) reg_16(
    .clk(reg_16__clk),
    .in(reg_16__in),
    .out(reg_16__out)
  );

  //Wire declarations for instance 'reg_17' (Module coreir_reg)
  wire  reg_17__clk;
  wire [15:0] reg_17__in;
  wire [15:0] reg_17__out;
  coreir_reg #(.clk_posedge(1),.init(16'bxxxxxxxxxxxxxxxx),.width(16)) reg_17(
    .clk(reg_17__clk),
    .in(reg_17__in),
    .out(reg_17__out)
  );

  //Wire declarations for instance 'reg_18' (Module coreir_reg)
  wire  reg_18__clk;
  wire [15:0] reg_18__in;
  wire [15:0] reg_18__out;
  coreir_reg #(.clk_posedge(1),.init(16'bxxxxxxxxxxxxxxxx),.width(16)) reg_18(
    .clk(reg_18__clk),
    .in(reg_18__in),
    .out(reg_18__out)
  );

  //Wire declarations for instance 'reg_19' (Module coreir_reg)
  wire  reg_19__clk;
  wire [15:0] reg_19__in;
  wire [15:0] reg_19__out;
  coreir_reg #(.clk_posedge(1),.init(16'bxxxxxxxxxxxxxxxx),.width(16)) reg_19(
    .clk(reg_19__clk),
    .in(reg_19__in),
    .out(reg_19__out)
  );

  //Wire declarations for instance 'reg_2' (Module coreir_reg)
  wire  reg_2__clk;
  wire [15:0] reg_2__in;
  wire [15:0] reg_2__out;
  coreir_reg #(.clk_posedge(1),.init(16'bxxxxxxxxxxxxxxxx),.width(16)) reg_2(
    .clk(reg_2__clk),
    .in(reg_2__in),
    .out(reg_2__out)
  );

  //Wire declarations for instance 'reg_3' (Module coreir_reg)
  wire  reg_3__clk;
  wire [15:0] reg_3__in;
  wire [15:0] reg_3__out;
  coreir_reg #(.clk_posedge(1),.init(16'bxxxxxxxxxxxxxxxx),.width(16)) reg_3(
    .clk(reg_3__clk),
    .in(reg_3__in),
    .out(reg_3__out)
  );

  //Wire declarations for instance 'reg_4' (Module coreir_reg)
  wire  reg_4__clk;
  wire [15:0] reg_4__in;
  wire [15:0] reg_4__out;
  coreir_reg #(.clk_posedge(1),.init(16'bxxxxxxxxxxxxxxxx),.width(16)) reg_4(
    .clk(reg_4__clk),
    .in(reg_4__in),
    .out(reg_4__out)
  );

  //Wire declarations for instance 'reg_5' (Module coreir_reg)
  wire  reg_5__clk;
  wire [15:0] reg_5__in;
  wire [15:0] reg_5__out;
  coreir_reg #(.clk_posedge(1),.init(16'bxxxxxxxxxxxxxxxx),.width(16)) reg_5(
    .clk(reg_5__clk),
    .in(reg_5__in),
    .out(reg_5__out)
  );

  //Wire declarations for instance 'reg_6' (Module coreir_reg)
  wire  reg_6__clk;
  wire [15:0] reg_6__in;
  wire [15:0] reg_6__out;
  coreir_reg #(.clk_posedge(1),.init(16'bxxxxxxxxxxxxxxxx),.width(16)) reg_6(
    .clk(reg_6__clk),
    .in(reg_6__in),
    .out(reg_6__out)
  );

  //Wire declarations for instance 'reg_7' (Module coreir_reg)
  wire  reg_7__clk;
  wire [15:0] reg_7__in;
  wire [15:0] reg_7__out;
  coreir_reg #(.clk_posedge(1),.init(16'bxxxxxxxxxxxxxxxx),.width(16)) reg_7(
    .clk(reg_7__clk),
    .in(reg_7__in),
    .out(reg_7__out)
  );

  //Wire declarations for instance 'reg_8' (Module coreir_reg)
  wire  reg_8__clk;
  wire [15:0] reg_8__in;
  wire [15:0] reg_8__out;
  coreir_reg #(.clk_posedge(1),.init(16'bxxxxxxxxxxxxxxxx),.width(16)) reg_8(
    .clk(reg_8__clk),
    .in(reg_8__in),
    .out(reg_8__out)
  );

  //Wire declarations for instance 'reg_9' (Module coreir_reg)
  wire  reg_9__clk;
  wire [15:0] reg_9__in;
  wire [15:0] reg_9__out;
  coreir_reg #(.clk_posedge(1),.init(16'bxxxxxxxxxxxxxxxx),.width(16)) reg_9(
    .clk(reg_9__clk),
    .in(reg_9__in),
    .out(reg_9__out)
  );

  //All the connections
  assign reg_1__in[15:0] = in_0[15:0];
  assign reg_2__in[15:0] = reg_1__out[15:0];
  assign out_18[15:0] = reg_1__out[15:0];
  assign reg_3__in[15:0] = reg_2__out[15:0];
  assign out_17[15:0] = reg_2__out[15:0];
  assign reg_4__in[15:0] = reg_3__out[15:0];
  assign out_16[15:0] = reg_3__out[15:0];
  assign reg_5__in[15:0] = reg_4__out[15:0];
  assign out_15[15:0] = reg_4__out[15:0];
  assign reg_6__in[15:0] = reg_5__out[15:0];
  assign out_14[15:0] = reg_5__out[15:0];
  assign reg_7__in[15:0] = reg_6__out[15:0];
  assign out_13[15:0] = reg_6__out[15:0];
  assign reg_8__in[15:0] = reg_7__out[15:0];
  assign out_12[15:0] = reg_7__out[15:0];
  assign reg_9__in[15:0] = reg_8__out[15:0];
  assign out_11[15:0] = reg_8__out[15:0];
  assign reg_10__in[15:0] = reg_9__out[15:0];
  assign out_10[15:0] = reg_9__out[15:0];
  assign reg_11__in[15:0] = reg_10__out[15:0];
  assign out_9[15:0] = reg_10__out[15:0];
  assign reg_12__in[15:0] = reg_11__out[15:0];
  assign out_8[15:0] = reg_11__out[15:0];
  assign reg_13__in[15:0] = reg_12__out[15:0];
  assign out_7[15:0] = reg_12__out[15:0];
  assign reg_14__in[15:0] = reg_13__out[15:0];
  assign out_6[15:0] = reg_13__out[15:0];
  assign reg_15__in[15:0] = reg_14__out[15:0];
  assign out_5[15:0] = reg_14__out[15:0];
  assign reg_16__in[15:0] = reg_15__out[15:0];
  assign out_4[15:0] = reg_15__out[15:0];
  assign reg_17__in[15:0] = reg_16__out[15:0];
  assign out_3[15:0] = reg_16__out[15:0];
  assign reg_18__in[15:0] = reg_17__out[15:0];
  assign out_2[15:0] = reg_17__out[15:0];
  assign reg_19__in[15:0] = reg_18__out[15:0];
  assign out_1[15:0] = reg_18__out[15:0];
  assign out_0[15:0] = reg_19__out[15:0];
  assign valid = wen;
  assign valid_chain = wen;
  assign reg_1__clk = clk;
  assign reg_12__clk = clk;
  assign reg_10__clk = clk;
  assign reg_11__clk = clk;
  assign reg_13__clk = clk;
  assign reg_14__clk = clk;
  assign reg_15__clk = clk;
  assign reg_16__clk = clk;
  assign reg_17__clk = clk;
  assign reg_18__clk = clk;
  assign reg_19__clk = clk;
  assign reg_2__clk = clk;
  assign reg_3__clk = clk;
  assign reg_4__clk = clk;
  assign reg_5__clk = clk;
  assign reg_6__clk = clk;
  assign reg_7__clk = clk;
  assign reg_8__clk = clk;
  assign reg_9__clk = clk;
  assign out_19[15:0] = in_0[15:0];

endmodule //linebuffer_U3

module reg_U25 #(parameter init=1) (
  input  clk,
  input  clr,
  input  en,
  input [8:0] in,
  output [8:0] out
);
  //Wire declarations for instance 'c0' (Module coreir_const)
  wire [8:0] c0__out;
  coreir_const #(.value(9'b000000000),.width(9)) c0(
    .out(c0__out)
  );

  //Wire declarations for instance 'clrMux' (Module coreir_mux)
  wire [8:0] clrMux__in0;
  wire [8:0] clrMux__in1;
  wire [8:0] clrMux__out;
  wire  clrMux__sel;
  coreir_mux #(.width(9)) clrMux(
    .in0(clrMux__in0),
    .in1(clrMux__in1),
    .out(clrMux__out),
    .sel(clrMux__sel)
  );

  //Wire declarations for instance 'enMux' (Module coreir_mux)
  wire [8:0] enMux__in0;
  wire [8:0] enMux__in1;
  wire [8:0] enMux__out;
  wire  enMux__sel;
  coreir_mux #(.width(9)) enMux(
    .in0(enMux__in0),
    .in1(enMux__in1),
    .out(enMux__out),
    .sel(enMux__sel)
  );

  //Wire declarations for instance 'reg0' (Module coreir_reg)
  wire  reg0__clk;
  wire [8:0] reg0__in;
  wire [8:0] reg0__out;
  coreir_reg #(.clk_posedge(1),.init(init),.width(9)) reg0(
    .clk(reg0__clk),
    .in(reg0__in),
    .out(reg0__out)
  );

  //All the connections
  assign reg0__in[8:0] = enMux__out[8:0];
  assign out[8:0] = reg0__out[8:0];
  assign enMux__in0[8:0] = reg0__out[8:0];
  assign reg0__clk = clk;
  assign enMux__sel = en;
  assign enMux__in1[8:0] = clrMux__out[8:0];
  assign clrMux__in1[8:0] = c0__out[8:0];
  assign clrMux__sel = clr;
  assign clrMux__in0[8:0] = in[8:0];

endmodule //reg_U25

module counter_U11 #(parameter init=1, parameter max=1) (
  input  clk,
  input  en,
  output [8:0] out,
  input  srst
);
  //Wire declarations for instance 'add' (Module coreir_add)
  wire [8:0] add__in0;
  wire [8:0] add__in1;
  wire [8:0] add__out;
  coreir_add #(.width(9)) add(
    .in0(add__in0),
    .in1(add__in1),
    .out(add__out)
  );

  //Wire declarations for instance 'c0' (Module coreir_const)
  wire [8:0] c0__out;
  coreir_const #(.value(9'b000000000),.width(9)) c0(
    .out(c0__out)
  );

  //Wire declarations for instance 'c1' (Module coreir_const)
  wire [8:0] c1__out;
  coreir_const #(.value(9'b000000001),.width(9)) c1(
    .out(c1__out)
  );

  //Wire declarations for instance 'eq' (Module coreir_eq)
  wire [8:0] eq__in0;
  wire [8:0] eq__in1;
  wire  eq__out;
  coreir_eq #(.width(9)) eq(
    .in0(eq__in0),
    .in1(eq__in1),
    .out(eq__out)
  );

  //Wire declarations for instance 'maxval' (Module coreir_const)
  wire [8:0] maxval__out;
  coreir_const #(.value(max),.width(9)) maxval(
    .out(maxval__out)
  );

  //Wire declarations for instance 'mux' (Module coreir_mux)
  wire [8:0] mux__in0;
  wire [8:0] mux__in1;
  wire [8:0] mux__out;
  wire  mux__sel;
  coreir_mux #(.width(9)) mux(
    .in0(mux__in0),
    .in1(mux__in1),
    .out(mux__out),
    .sel(mux__sel)
  );

  //Wire declarations for instance 'r' (Module reg_U25)
  wire  r__clk;
  wire  r__clr;
  wire  r__en;
  wire [8:0] r__in;
  wire [8:0] r__out;
  reg_U25 #(.init(init)) r(
    .clk(r__clk),
    .clr(r__clr),
    .en(r__en),
    .in(r__in),
    .out(r__out)
  );

  //All the connections
  assign r__clk = clk;
  assign r__en = en;
  assign r__clr = srst;
  assign add__in1[8:0] = c1__out[8:0];
  assign add__in0[8:0] = r__out[8:0];
  assign out[8:0] = r__out[8:0];
  assign eq__in0[8:0] = r__out[8:0];
  assign mux__sel = eq__out;
  assign eq__in1[8:0] = maxval__out[8:0];
  assign mux__in0[8:0] = add__out[8:0];
  assign mux__in1[8:0] = c0__out[8:0];
  assign r__in[8:0] = mux__out[8:0];

endmodule //counter_U11

module coreir_ule #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output out
);
  assign out = in0 <= in1;

endmodule //coreir_ule

module coreir_ult #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output out
);
  assign out = in0 < in1;

endmodule //coreir_ult

module coreir_const160 (
  output [15:0] out
);
  //Wire declarations for instance 'bit_const_GND' (Module corebit_const)
  wire  bit_const_GND__out;
  corebit_const #(.value(0)) bit_const_GND(
    .out(bit_const_GND__out)
  );

  //All the connections
  assign out[0] = bit_const_GND__out;
  assign out[11] = bit_const_GND__out;
  assign out[12] = bit_const_GND__out;
  assign out[13] = bit_const_GND__out;
  assign out[14] = bit_const_GND__out;
  assign out[15] = bit_const_GND__out;
  assign out[1] = bit_const_GND__out;
  assign out[2] = bit_const_GND__out;
  assign out[3] = bit_const_GND__out;
  assign out[4] = bit_const_GND__out;
  assign out[5] = bit_const_GND__out;
  assign out[6] = bit_const_GND__out;
  assign out[7] = bit_const_GND__out;
  assign out[8] = bit_const_GND__out;
  assign out[10] = bit_const_GND__out;
  assign out[9] = bit_const_GND__out;

endmodule //coreir_const160

module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ (
  input [15:0] in0,
  input [15:0] in1,
  output [15:0] out
);
  //Wire declarations for instance 'inst0' (Module Add16)
  wire [15:0] inst0__I0;
  wire [15:0] inst0__I1;
  wire [15:0] inst0__O;
  Add16 inst0(
    .I0(inst0__I0),
    .I1(inst0__I1),
    .O(inst0__O)
  );

  //All the connections
  assign inst0__I0[15:0] = in0[15:0];
  assign inst0__I1[15:0] = in1[15:0];
  assign out[15:0] = inst0__O[15:0];

endmodule //renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___

module reduceParallelPower2Inputs_U2 (
  input [15:0] in_0,
  input [15:0] in_1,
  input [15:0] in_10,
  input [15:0] in_100,
  input [15:0] in_101,
  input [15:0] in_102,
  input [15:0] in_103,
  input [15:0] in_104,
  input [15:0] in_105,
  input [15:0] in_106,
  input [15:0] in_107,
  input [15:0] in_108,
  input [15:0] in_109,
  input [15:0] in_11,
  input [15:0] in_110,
  input [15:0] in_111,
  input [15:0] in_112,
  input [15:0] in_113,
  input [15:0] in_114,
  input [15:0] in_115,
  input [15:0] in_116,
  input [15:0] in_117,
  input [15:0] in_118,
  input [15:0] in_119,
  input [15:0] in_12,
  input [15:0] in_120,
  input [15:0] in_121,
  input [15:0] in_122,
  input [15:0] in_123,
  input [15:0] in_124,
  input [15:0] in_125,
  input [15:0] in_126,
  input [15:0] in_127,
  input [15:0] in_128,
  input [15:0] in_129,
  input [15:0] in_13,
  input [15:0] in_130,
  input [15:0] in_131,
  input [15:0] in_132,
  input [15:0] in_133,
  input [15:0] in_134,
  input [15:0] in_135,
  input [15:0] in_136,
  input [15:0] in_137,
  input [15:0] in_138,
  input [15:0] in_139,
  input [15:0] in_14,
  input [15:0] in_140,
  input [15:0] in_141,
  input [15:0] in_142,
  input [15:0] in_143,
  input [15:0] in_144,
  input [15:0] in_145,
  input [15:0] in_146,
  input [15:0] in_147,
  input [15:0] in_148,
  input [15:0] in_149,
  input [15:0] in_15,
  input [15:0] in_150,
  input [15:0] in_151,
  input [15:0] in_152,
  input [15:0] in_153,
  input [15:0] in_154,
  input [15:0] in_155,
  input [15:0] in_156,
  input [15:0] in_157,
  input [15:0] in_158,
  input [15:0] in_159,
  input [15:0] in_16,
  input [15:0] in_160,
  input [15:0] in_161,
  input [15:0] in_162,
  input [15:0] in_163,
  input [15:0] in_164,
  input [15:0] in_165,
  input [15:0] in_166,
  input [15:0] in_167,
  input [15:0] in_168,
  input [15:0] in_169,
  input [15:0] in_17,
  input [15:0] in_170,
  input [15:0] in_171,
  input [15:0] in_172,
  input [15:0] in_173,
  input [15:0] in_174,
  input [15:0] in_175,
  input [15:0] in_176,
  input [15:0] in_177,
  input [15:0] in_178,
  input [15:0] in_179,
  input [15:0] in_18,
  input [15:0] in_180,
  input [15:0] in_181,
  input [15:0] in_182,
  input [15:0] in_183,
  input [15:0] in_184,
  input [15:0] in_185,
  input [15:0] in_186,
  input [15:0] in_187,
  input [15:0] in_188,
  input [15:0] in_189,
  input [15:0] in_19,
  input [15:0] in_190,
  input [15:0] in_191,
  input [15:0] in_192,
  input [15:0] in_193,
  input [15:0] in_194,
  input [15:0] in_195,
  input [15:0] in_196,
  input [15:0] in_197,
  input [15:0] in_198,
  input [15:0] in_199,
  input [15:0] in_2,
  input [15:0] in_20,
  input [15:0] in_200,
  input [15:0] in_201,
  input [15:0] in_202,
  input [15:0] in_203,
  input [15:0] in_204,
  input [15:0] in_205,
  input [15:0] in_206,
  input [15:0] in_207,
  input [15:0] in_208,
  input [15:0] in_209,
  input [15:0] in_21,
  input [15:0] in_210,
  input [15:0] in_211,
  input [15:0] in_212,
  input [15:0] in_213,
  input [15:0] in_214,
  input [15:0] in_215,
  input [15:0] in_216,
  input [15:0] in_217,
  input [15:0] in_218,
  input [15:0] in_219,
  input [15:0] in_22,
  input [15:0] in_220,
  input [15:0] in_221,
  input [15:0] in_222,
  input [15:0] in_223,
  input [15:0] in_224,
  input [15:0] in_225,
  input [15:0] in_226,
  input [15:0] in_227,
  input [15:0] in_228,
  input [15:0] in_229,
  input [15:0] in_23,
  input [15:0] in_230,
  input [15:0] in_231,
  input [15:0] in_232,
  input [15:0] in_233,
  input [15:0] in_234,
  input [15:0] in_235,
  input [15:0] in_236,
  input [15:0] in_237,
  input [15:0] in_238,
  input [15:0] in_239,
  input [15:0] in_24,
  input [15:0] in_240,
  input [15:0] in_241,
  input [15:0] in_242,
  input [15:0] in_243,
  input [15:0] in_244,
  input [15:0] in_245,
  input [15:0] in_246,
  input [15:0] in_247,
  input [15:0] in_248,
  input [15:0] in_249,
  input [15:0] in_25,
  input [15:0] in_250,
  input [15:0] in_251,
  input [15:0] in_252,
  input [15:0] in_253,
  input [15:0] in_254,
  input [15:0] in_255,
  input [15:0] in_256,
  input [15:0] in_257,
  input [15:0] in_258,
  input [15:0] in_259,
  input [15:0] in_26,
  input [15:0] in_260,
  input [15:0] in_261,
  input [15:0] in_262,
  input [15:0] in_263,
  input [15:0] in_264,
  input [15:0] in_265,
  input [15:0] in_266,
  input [15:0] in_267,
  input [15:0] in_268,
  input [15:0] in_269,
  input [15:0] in_27,
  input [15:0] in_270,
  input [15:0] in_271,
  input [15:0] in_272,
  input [15:0] in_273,
  input [15:0] in_274,
  input [15:0] in_275,
  input [15:0] in_276,
  input [15:0] in_277,
  input [15:0] in_278,
  input [15:0] in_279,
  input [15:0] in_28,
  input [15:0] in_280,
  input [15:0] in_281,
  input [15:0] in_282,
  input [15:0] in_283,
  input [15:0] in_284,
  input [15:0] in_285,
  input [15:0] in_286,
  input [15:0] in_287,
  input [15:0] in_288,
  input [15:0] in_289,
  input [15:0] in_29,
  input [15:0] in_290,
  input [15:0] in_291,
  input [15:0] in_292,
  input [15:0] in_293,
  input [15:0] in_294,
  input [15:0] in_295,
  input [15:0] in_296,
  input [15:0] in_297,
  input [15:0] in_298,
  input [15:0] in_299,
  input [15:0] in_3,
  input [15:0] in_30,
  input [15:0] in_300,
  input [15:0] in_301,
  input [15:0] in_302,
  input [15:0] in_303,
  input [15:0] in_304,
  input [15:0] in_305,
  input [15:0] in_306,
  input [15:0] in_307,
  input [15:0] in_308,
  input [15:0] in_309,
  input [15:0] in_31,
  input [15:0] in_310,
  input [15:0] in_311,
  input [15:0] in_312,
  input [15:0] in_313,
  input [15:0] in_314,
  input [15:0] in_315,
  input [15:0] in_316,
  input [15:0] in_317,
  input [15:0] in_318,
  input [15:0] in_319,
  input [15:0] in_32,
  input [15:0] in_320,
  input [15:0] in_321,
  input [15:0] in_322,
  input [15:0] in_323,
  input [15:0] in_324,
  input [15:0] in_325,
  input [15:0] in_326,
  input [15:0] in_327,
  input [15:0] in_328,
  input [15:0] in_329,
  input [15:0] in_33,
  input [15:0] in_330,
  input [15:0] in_331,
  input [15:0] in_332,
  input [15:0] in_333,
  input [15:0] in_334,
  input [15:0] in_335,
  input [15:0] in_336,
  input [15:0] in_337,
  input [15:0] in_338,
  input [15:0] in_339,
  input [15:0] in_34,
  input [15:0] in_340,
  input [15:0] in_341,
  input [15:0] in_342,
  input [15:0] in_343,
  input [15:0] in_344,
  input [15:0] in_345,
  input [15:0] in_346,
  input [15:0] in_347,
  input [15:0] in_348,
  input [15:0] in_349,
  input [15:0] in_35,
  input [15:0] in_350,
  input [15:0] in_351,
  input [15:0] in_352,
  input [15:0] in_353,
  input [15:0] in_354,
  input [15:0] in_355,
  input [15:0] in_356,
  input [15:0] in_357,
  input [15:0] in_358,
  input [15:0] in_359,
  input [15:0] in_36,
  input [15:0] in_360,
  input [15:0] in_361,
  input [15:0] in_362,
  input [15:0] in_363,
  input [15:0] in_364,
  input [15:0] in_365,
  input [15:0] in_366,
  input [15:0] in_367,
  input [15:0] in_368,
  input [15:0] in_369,
  input [15:0] in_37,
  input [15:0] in_370,
  input [15:0] in_371,
  input [15:0] in_372,
  input [15:0] in_373,
  input [15:0] in_374,
  input [15:0] in_375,
  input [15:0] in_376,
  input [15:0] in_377,
  input [15:0] in_378,
  input [15:0] in_379,
  input [15:0] in_38,
  input [15:0] in_380,
  input [15:0] in_381,
  input [15:0] in_382,
  input [15:0] in_383,
  input [15:0] in_384,
  input [15:0] in_385,
  input [15:0] in_386,
  input [15:0] in_387,
  input [15:0] in_388,
  input [15:0] in_389,
  input [15:0] in_39,
  input [15:0] in_390,
  input [15:0] in_391,
  input [15:0] in_392,
  input [15:0] in_393,
  input [15:0] in_394,
  input [15:0] in_395,
  input [15:0] in_396,
  input [15:0] in_397,
  input [15:0] in_398,
  input [15:0] in_399,
  input [15:0] in_4,
  input [15:0] in_40,
  input [15:0] in_400,
  input [15:0] in_401,
  input [15:0] in_402,
  input [15:0] in_403,
  input [15:0] in_404,
  input [15:0] in_405,
  input [15:0] in_406,
  input [15:0] in_407,
  input [15:0] in_408,
  input [15:0] in_409,
  input [15:0] in_41,
  input [15:0] in_410,
  input [15:0] in_411,
  input [15:0] in_412,
  input [15:0] in_413,
  input [15:0] in_414,
  input [15:0] in_415,
  input [15:0] in_416,
  input [15:0] in_417,
  input [15:0] in_418,
  input [15:0] in_419,
  input [15:0] in_42,
  input [15:0] in_420,
  input [15:0] in_421,
  input [15:0] in_422,
  input [15:0] in_423,
  input [15:0] in_424,
  input [15:0] in_425,
  input [15:0] in_426,
  input [15:0] in_427,
  input [15:0] in_428,
  input [15:0] in_429,
  input [15:0] in_43,
  input [15:0] in_430,
  input [15:0] in_431,
  input [15:0] in_432,
  input [15:0] in_433,
  input [15:0] in_434,
  input [15:0] in_435,
  input [15:0] in_436,
  input [15:0] in_437,
  input [15:0] in_438,
  input [15:0] in_439,
  input [15:0] in_44,
  input [15:0] in_440,
  input [15:0] in_441,
  input [15:0] in_442,
  input [15:0] in_443,
  input [15:0] in_444,
  input [15:0] in_445,
  input [15:0] in_446,
  input [15:0] in_447,
  input [15:0] in_448,
  input [15:0] in_449,
  input [15:0] in_45,
  input [15:0] in_450,
  input [15:0] in_451,
  input [15:0] in_452,
  input [15:0] in_453,
  input [15:0] in_454,
  input [15:0] in_455,
  input [15:0] in_456,
  input [15:0] in_457,
  input [15:0] in_458,
  input [15:0] in_459,
  input [15:0] in_46,
  input [15:0] in_460,
  input [15:0] in_461,
  input [15:0] in_462,
  input [15:0] in_463,
  input [15:0] in_464,
  input [15:0] in_465,
  input [15:0] in_466,
  input [15:0] in_467,
  input [15:0] in_468,
  input [15:0] in_469,
  input [15:0] in_47,
  input [15:0] in_470,
  input [15:0] in_471,
  input [15:0] in_472,
  input [15:0] in_473,
  input [15:0] in_474,
  input [15:0] in_475,
  input [15:0] in_476,
  input [15:0] in_477,
  input [15:0] in_478,
  input [15:0] in_479,
  input [15:0] in_48,
  input [15:0] in_480,
  input [15:0] in_481,
  input [15:0] in_482,
  input [15:0] in_483,
  input [15:0] in_484,
  input [15:0] in_485,
  input [15:0] in_486,
  input [15:0] in_487,
  input [15:0] in_488,
  input [15:0] in_489,
  input [15:0] in_49,
  input [15:0] in_490,
  input [15:0] in_491,
  input [15:0] in_492,
  input [15:0] in_493,
  input [15:0] in_494,
  input [15:0] in_495,
  input [15:0] in_496,
  input [15:0] in_497,
  input [15:0] in_498,
  input [15:0] in_499,
  input [15:0] in_5,
  input [15:0] in_50,
  input [15:0] in_500,
  input [15:0] in_501,
  input [15:0] in_502,
  input [15:0] in_503,
  input [15:0] in_504,
  input [15:0] in_505,
  input [15:0] in_506,
  input [15:0] in_507,
  input [15:0] in_508,
  input [15:0] in_509,
  input [15:0] in_51,
  input [15:0] in_510,
  input [15:0] in_511,
  input [15:0] in_52,
  input [15:0] in_53,
  input [15:0] in_54,
  input [15:0] in_55,
  input [15:0] in_56,
  input [15:0] in_57,
  input [15:0] in_58,
  input [15:0] in_59,
  input [15:0] in_6,
  input [15:0] in_60,
  input [15:0] in_61,
  input [15:0] in_62,
  input [15:0] in_63,
  input [15:0] in_64,
  input [15:0] in_65,
  input [15:0] in_66,
  input [15:0] in_67,
  input [15:0] in_68,
  input [15:0] in_69,
  input [15:0] in_7,
  input [15:0] in_70,
  input [15:0] in_71,
  input [15:0] in_72,
  input [15:0] in_73,
  input [15:0] in_74,
  input [15:0] in_75,
  input [15:0] in_76,
  input [15:0] in_77,
  input [15:0] in_78,
  input [15:0] in_79,
  input [15:0] in_8,
  input [15:0] in_80,
  input [15:0] in_81,
  input [15:0] in_82,
  input [15:0] in_83,
  input [15:0] in_84,
  input [15:0] in_85,
  input [15:0] in_86,
  input [15:0] in_87,
  input [15:0] in_88,
  input [15:0] in_89,
  input [15:0] in_9,
  input [15:0] in_90,
  input [15:0] in_91,
  input [15:0] in_92,
  input [15:0] in_93,
  input [15:0] in_94,
  input [15:0] in_95,
  input [15:0] in_96,
  input [15:0] in_97,
  input [15:0] in_98,
  input [15:0] in_99,
  output [15:0] out
);
  //Wire declarations for instance 'op_0_0' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_0_0__in0;
  wire [15:0] op_0_0__in1;
  wire [15:0] op_0_0__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_0_0(
    .in0(op_0_0__in0),
    .in1(op_0_0__in1),
    .out(op_0_0__out)
  );

  //Wire declarations for instance 'op_1_0' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_1_0__in0;
  wire [15:0] op_1_0__in1;
  wire [15:0] op_1_0__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_1_0(
    .in0(op_1_0__in0),
    .in1(op_1_0__in1),
    .out(op_1_0__out)
  );

  //Wire declarations for instance 'op_1_1' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_1_1__in0;
  wire [15:0] op_1_1__in1;
  wire [15:0] op_1_1__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_1_1(
    .in0(op_1_1__in0),
    .in1(op_1_1__in1),
    .out(op_1_1__out)
  );

  //Wire declarations for instance 'op_2_0' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_2_0__in0;
  wire [15:0] op_2_0__in1;
  wire [15:0] op_2_0__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_2_0(
    .in0(op_2_0__in0),
    .in1(op_2_0__in1),
    .out(op_2_0__out)
  );

  //Wire declarations for instance 'op_2_1' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_2_1__in0;
  wire [15:0] op_2_1__in1;
  wire [15:0] op_2_1__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_2_1(
    .in0(op_2_1__in0),
    .in1(op_2_1__in1),
    .out(op_2_1__out)
  );

  //Wire declarations for instance 'op_2_2' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_2_2__in0;
  wire [15:0] op_2_2__in1;
  wire [15:0] op_2_2__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_2_2(
    .in0(op_2_2__in0),
    .in1(op_2_2__in1),
    .out(op_2_2__out)
  );

  //Wire declarations for instance 'op_2_3' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_2_3__in0;
  wire [15:0] op_2_3__in1;
  wire [15:0] op_2_3__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_2_3(
    .in0(op_2_3__in0),
    .in1(op_2_3__in1),
    .out(op_2_3__out)
  );

  //Wire declarations for instance 'op_3_0' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_3_0__in0;
  wire [15:0] op_3_0__in1;
  wire [15:0] op_3_0__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_3_0(
    .in0(op_3_0__in0),
    .in1(op_3_0__in1),
    .out(op_3_0__out)
  );

  //Wire declarations for instance 'op_3_1' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_3_1__in0;
  wire [15:0] op_3_1__in1;
  wire [15:0] op_3_1__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_3_1(
    .in0(op_3_1__in0),
    .in1(op_3_1__in1),
    .out(op_3_1__out)
  );

  //Wire declarations for instance 'op_3_2' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_3_2__in0;
  wire [15:0] op_3_2__in1;
  wire [15:0] op_3_2__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_3_2(
    .in0(op_3_2__in0),
    .in1(op_3_2__in1),
    .out(op_3_2__out)
  );

  //Wire declarations for instance 'op_3_3' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_3_3__in0;
  wire [15:0] op_3_3__in1;
  wire [15:0] op_3_3__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_3_3(
    .in0(op_3_3__in0),
    .in1(op_3_3__in1),
    .out(op_3_3__out)
  );

  //Wire declarations for instance 'op_3_4' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_3_4__in0;
  wire [15:0] op_3_4__in1;
  wire [15:0] op_3_4__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_3_4(
    .in0(op_3_4__in0),
    .in1(op_3_4__in1),
    .out(op_3_4__out)
  );

  //Wire declarations for instance 'op_3_5' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_3_5__in0;
  wire [15:0] op_3_5__in1;
  wire [15:0] op_3_5__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_3_5(
    .in0(op_3_5__in0),
    .in1(op_3_5__in1),
    .out(op_3_5__out)
  );

  //Wire declarations for instance 'op_3_6' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_3_6__in0;
  wire [15:0] op_3_6__in1;
  wire [15:0] op_3_6__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_3_6(
    .in0(op_3_6__in0),
    .in1(op_3_6__in1),
    .out(op_3_6__out)
  );

  //Wire declarations for instance 'op_3_7' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_3_7__in0;
  wire [15:0] op_3_7__in1;
  wire [15:0] op_3_7__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_3_7(
    .in0(op_3_7__in0),
    .in1(op_3_7__in1),
    .out(op_3_7__out)
  );

  //Wire declarations for instance 'op_4_0' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_4_0__in0;
  wire [15:0] op_4_0__in1;
  wire [15:0] op_4_0__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_4_0(
    .in0(op_4_0__in0),
    .in1(op_4_0__in1),
    .out(op_4_0__out)
  );

  //Wire declarations for instance 'op_4_1' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_4_1__in0;
  wire [15:0] op_4_1__in1;
  wire [15:0] op_4_1__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_4_1(
    .in0(op_4_1__in0),
    .in1(op_4_1__in1),
    .out(op_4_1__out)
  );

  //Wire declarations for instance 'op_4_10' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_4_10__in0;
  wire [15:0] op_4_10__in1;
  wire [15:0] op_4_10__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_4_10(
    .in0(op_4_10__in0),
    .in1(op_4_10__in1),
    .out(op_4_10__out)
  );

  //Wire declarations for instance 'op_4_11' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_4_11__in0;
  wire [15:0] op_4_11__in1;
  wire [15:0] op_4_11__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_4_11(
    .in0(op_4_11__in0),
    .in1(op_4_11__in1),
    .out(op_4_11__out)
  );

  //Wire declarations for instance 'op_4_12' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_4_12__in0;
  wire [15:0] op_4_12__in1;
  wire [15:0] op_4_12__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_4_12(
    .in0(op_4_12__in0),
    .in1(op_4_12__in1),
    .out(op_4_12__out)
  );

  //Wire declarations for instance 'op_4_13' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_4_13__in0;
  wire [15:0] op_4_13__in1;
  wire [15:0] op_4_13__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_4_13(
    .in0(op_4_13__in0),
    .in1(op_4_13__in1),
    .out(op_4_13__out)
  );

  //Wire declarations for instance 'op_4_14' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_4_14__in0;
  wire [15:0] op_4_14__in1;
  wire [15:0] op_4_14__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_4_14(
    .in0(op_4_14__in0),
    .in1(op_4_14__in1),
    .out(op_4_14__out)
  );

  //Wire declarations for instance 'op_4_15' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_4_15__in0;
  wire [15:0] op_4_15__in1;
  wire [15:0] op_4_15__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_4_15(
    .in0(op_4_15__in0),
    .in1(op_4_15__in1),
    .out(op_4_15__out)
  );

  //Wire declarations for instance 'op_4_2' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_4_2__in0;
  wire [15:0] op_4_2__in1;
  wire [15:0] op_4_2__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_4_2(
    .in0(op_4_2__in0),
    .in1(op_4_2__in1),
    .out(op_4_2__out)
  );

  //Wire declarations for instance 'op_4_3' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_4_3__in0;
  wire [15:0] op_4_3__in1;
  wire [15:0] op_4_3__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_4_3(
    .in0(op_4_3__in0),
    .in1(op_4_3__in1),
    .out(op_4_3__out)
  );

  //Wire declarations for instance 'op_4_4' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_4_4__in0;
  wire [15:0] op_4_4__in1;
  wire [15:0] op_4_4__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_4_4(
    .in0(op_4_4__in0),
    .in1(op_4_4__in1),
    .out(op_4_4__out)
  );

  //Wire declarations for instance 'op_4_5' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_4_5__in0;
  wire [15:0] op_4_5__in1;
  wire [15:0] op_4_5__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_4_5(
    .in0(op_4_5__in0),
    .in1(op_4_5__in1),
    .out(op_4_5__out)
  );

  //Wire declarations for instance 'op_4_6' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_4_6__in0;
  wire [15:0] op_4_6__in1;
  wire [15:0] op_4_6__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_4_6(
    .in0(op_4_6__in0),
    .in1(op_4_6__in1),
    .out(op_4_6__out)
  );

  //Wire declarations for instance 'op_4_7' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_4_7__in0;
  wire [15:0] op_4_7__in1;
  wire [15:0] op_4_7__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_4_7(
    .in0(op_4_7__in0),
    .in1(op_4_7__in1),
    .out(op_4_7__out)
  );

  //Wire declarations for instance 'op_4_8' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_4_8__in0;
  wire [15:0] op_4_8__in1;
  wire [15:0] op_4_8__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_4_8(
    .in0(op_4_8__in0),
    .in1(op_4_8__in1),
    .out(op_4_8__out)
  );

  //Wire declarations for instance 'op_4_9' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_4_9__in0;
  wire [15:0] op_4_9__in1;
  wire [15:0] op_4_9__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_4_9(
    .in0(op_4_9__in0),
    .in1(op_4_9__in1),
    .out(op_4_9__out)
  );

  //Wire declarations for instance 'op_5_0' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_0__in0;
  wire [15:0] op_5_0__in1;
  wire [15:0] op_5_0__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_0(
    .in0(op_5_0__in0),
    .in1(op_5_0__in1),
    .out(op_5_0__out)
  );

  //Wire declarations for instance 'op_5_1' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_1__in0;
  wire [15:0] op_5_1__in1;
  wire [15:0] op_5_1__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_1(
    .in0(op_5_1__in0),
    .in1(op_5_1__in1),
    .out(op_5_1__out)
  );

  //Wire declarations for instance 'op_5_10' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_10__in0;
  wire [15:0] op_5_10__in1;
  wire [15:0] op_5_10__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_10(
    .in0(op_5_10__in0),
    .in1(op_5_10__in1),
    .out(op_5_10__out)
  );

  //Wire declarations for instance 'op_5_11' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_11__in0;
  wire [15:0] op_5_11__in1;
  wire [15:0] op_5_11__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_11(
    .in0(op_5_11__in0),
    .in1(op_5_11__in1),
    .out(op_5_11__out)
  );

  //Wire declarations for instance 'op_5_12' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_12__in0;
  wire [15:0] op_5_12__in1;
  wire [15:0] op_5_12__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_12(
    .in0(op_5_12__in0),
    .in1(op_5_12__in1),
    .out(op_5_12__out)
  );

  //Wire declarations for instance 'op_5_13' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_13__in0;
  wire [15:0] op_5_13__in1;
  wire [15:0] op_5_13__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_13(
    .in0(op_5_13__in0),
    .in1(op_5_13__in1),
    .out(op_5_13__out)
  );

  //Wire declarations for instance 'op_5_14' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_14__in0;
  wire [15:0] op_5_14__in1;
  wire [15:0] op_5_14__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_14(
    .in0(op_5_14__in0),
    .in1(op_5_14__in1),
    .out(op_5_14__out)
  );

  //Wire declarations for instance 'op_5_15' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_15__in0;
  wire [15:0] op_5_15__in1;
  wire [15:0] op_5_15__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_15(
    .in0(op_5_15__in0),
    .in1(op_5_15__in1),
    .out(op_5_15__out)
  );

  //Wire declarations for instance 'op_5_16' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_16__in0;
  wire [15:0] op_5_16__in1;
  wire [15:0] op_5_16__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_16(
    .in0(op_5_16__in0),
    .in1(op_5_16__in1),
    .out(op_5_16__out)
  );

  //Wire declarations for instance 'op_5_17' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_17__in0;
  wire [15:0] op_5_17__in1;
  wire [15:0] op_5_17__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_17(
    .in0(op_5_17__in0),
    .in1(op_5_17__in1),
    .out(op_5_17__out)
  );

  //Wire declarations for instance 'op_5_18' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_18__in0;
  wire [15:0] op_5_18__in1;
  wire [15:0] op_5_18__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_18(
    .in0(op_5_18__in0),
    .in1(op_5_18__in1),
    .out(op_5_18__out)
  );

  //Wire declarations for instance 'op_5_19' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_19__in0;
  wire [15:0] op_5_19__in1;
  wire [15:0] op_5_19__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_19(
    .in0(op_5_19__in0),
    .in1(op_5_19__in1),
    .out(op_5_19__out)
  );

  //Wire declarations for instance 'op_5_2' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_2__in0;
  wire [15:0] op_5_2__in1;
  wire [15:0] op_5_2__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_2(
    .in0(op_5_2__in0),
    .in1(op_5_2__in1),
    .out(op_5_2__out)
  );

  //Wire declarations for instance 'op_5_20' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_20__in0;
  wire [15:0] op_5_20__in1;
  wire [15:0] op_5_20__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_20(
    .in0(op_5_20__in0),
    .in1(op_5_20__in1),
    .out(op_5_20__out)
  );

  //Wire declarations for instance 'op_5_21' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_21__in0;
  wire [15:0] op_5_21__in1;
  wire [15:0] op_5_21__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_21(
    .in0(op_5_21__in0),
    .in1(op_5_21__in1),
    .out(op_5_21__out)
  );

  //Wire declarations for instance 'op_5_22' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_22__in0;
  wire [15:0] op_5_22__in1;
  wire [15:0] op_5_22__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_22(
    .in0(op_5_22__in0),
    .in1(op_5_22__in1),
    .out(op_5_22__out)
  );

  //Wire declarations for instance 'op_5_23' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_23__in0;
  wire [15:0] op_5_23__in1;
  wire [15:0] op_5_23__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_23(
    .in0(op_5_23__in0),
    .in1(op_5_23__in1),
    .out(op_5_23__out)
  );

  //Wire declarations for instance 'op_5_24' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_24__in0;
  wire [15:0] op_5_24__in1;
  wire [15:0] op_5_24__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_24(
    .in0(op_5_24__in0),
    .in1(op_5_24__in1),
    .out(op_5_24__out)
  );

  //Wire declarations for instance 'op_5_25' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_25__in0;
  wire [15:0] op_5_25__in1;
  wire [15:0] op_5_25__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_25(
    .in0(op_5_25__in0),
    .in1(op_5_25__in1),
    .out(op_5_25__out)
  );

  //Wire declarations for instance 'op_5_26' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_26__in0;
  wire [15:0] op_5_26__in1;
  wire [15:0] op_5_26__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_26(
    .in0(op_5_26__in0),
    .in1(op_5_26__in1),
    .out(op_5_26__out)
  );

  //Wire declarations for instance 'op_5_27' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_27__in0;
  wire [15:0] op_5_27__in1;
  wire [15:0] op_5_27__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_27(
    .in0(op_5_27__in0),
    .in1(op_5_27__in1),
    .out(op_5_27__out)
  );

  //Wire declarations for instance 'op_5_28' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_28__in0;
  wire [15:0] op_5_28__in1;
  wire [15:0] op_5_28__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_28(
    .in0(op_5_28__in0),
    .in1(op_5_28__in1),
    .out(op_5_28__out)
  );

  //Wire declarations for instance 'op_5_29' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_29__in0;
  wire [15:0] op_5_29__in1;
  wire [15:0] op_5_29__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_29(
    .in0(op_5_29__in0),
    .in1(op_5_29__in1),
    .out(op_5_29__out)
  );

  //Wire declarations for instance 'op_5_3' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_3__in0;
  wire [15:0] op_5_3__in1;
  wire [15:0] op_5_3__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_3(
    .in0(op_5_3__in0),
    .in1(op_5_3__in1),
    .out(op_5_3__out)
  );

  //Wire declarations for instance 'op_5_30' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_30__in0;
  wire [15:0] op_5_30__in1;
  wire [15:0] op_5_30__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_30(
    .in0(op_5_30__in0),
    .in1(op_5_30__in1),
    .out(op_5_30__out)
  );

  //Wire declarations for instance 'op_5_31' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_31__in0;
  wire [15:0] op_5_31__in1;
  wire [15:0] op_5_31__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_31(
    .in0(op_5_31__in0),
    .in1(op_5_31__in1),
    .out(op_5_31__out)
  );

  //Wire declarations for instance 'op_5_4' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_4__in0;
  wire [15:0] op_5_4__in1;
  wire [15:0] op_5_4__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_4(
    .in0(op_5_4__in0),
    .in1(op_5_4__in1),
    .out(op_5_4__out)
  );

  //Wire declarations for instance 'op_5_5' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_5__in0;
  wire [15:0] op_5_5__in1;
  wire [15:0] op_5_5__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_5(
    .in0(op_5_5__in0),
    .in1(op_5_5__in1),
    .out(op_5_5__out)
  );

  //Wire declarations for instance 'op_5_6' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_6__in0;
  wire [15:0] op_5_6__in1;
  wire [15:0] op_5_6__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_6(
    .in0(op_5_6__in0),
    .in1(op_5_6__in1),
    .out(op_5_6__out)
  );

  //Wire declarations for instance 'op_5_7' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_7__in0;
  wire [15:0] op_5_7__in1;
  wire [15:0] op_5_7__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_7(
    .in0(op_5_7__in0),
    .in1(op_5_7__in1),
    .out(op_5_7__out)
  );

  //Wire declarations for instance 'op_5_8' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_8__in0;
  wire [15:0] op_5_8__in1;
  wire [15:0] op_5_8__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_8(
    .in0(op_5_8__in0),
    .in1(op_5_8__in1),
    .out(op_5_8__out)
  );

  //Wire declarations for instance 'op_5_9' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_5_9__in0;
  wire [15:0] op_5_9__in1;
  wire [15:0] op_5_9__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_5_9(
    .in0(op_5_9__in0),
    .in1(op_5_9__in1),
    .out(op_5_9__out)
  );

  //Wire declarations for instance 'op_6_0' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_0__in0;
  wire [15:0] op_6_0__in1;
  wire [15:0] op_6_0__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_0(
    .in0(op_6_0__in0),
    .in1(op_6_0__in1),
    .out(op_6_0__out)
  );

  //Wire declarations for instance 'op_6_1' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_1__in0;
  wire [15:0] op_6_1__in1;
  wire [15:0] op_6_1__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_1(
    .in0(op_6_1__in0),
    .in1(op_6_1__in1),
    .out(op_6_1__out)
  );

  //Wire declarations for instance 'op_6_10' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_10__in0;
  wire [15:0] op_6_10__in1;
  wire [15:0] op_6_10__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_10(
    .in0(op_6_10__in0),
    .in1(op_6_10__in1),
    .out(op_6_10__out)
  );

  //Wire declarations for instance 'op_6_11' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_11__in0;
  wire [15:0] op_6_11__in1;
  wire [15:0] op_6_11__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_11(
    .in0(op_6_11__in0),
    .in1(op_6_11__in1),
    .out(op_6_11__out)
  );

  //Wire declarations for instance 'op_6_12' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_12__in0;
  wire [15:0] op_6_12__in1;
  wire [15:0] op_6_12__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_12(
    .in0(op_6_12__in0),
    .in1(op_6_12__in1),
    .out(op_6_12__out)
  );

  //Wire declarations for instance 'op_6_13' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_13__in0;
  wire [15:0] op_6_13__in1;
  wire [15:0] op_6_13__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_13(
    .in0(op_6_13__in0),
    .in1(op_6_13__in1),
    .out(op_6_13__out)
  );

  //Wire declarations for instance 'op_6_14' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_14__in0;
  wire [15:0] op_6_14__in1;
  wire [15:0] op_6_14__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_14(
    .in0(op_6_14__in0),
    .in1(op_6_14__in1),
    .out(op_6_14__out)
  );

  //Wire declarations for instance 'op_6_15' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_15__in0;
  wire [15:0] op_6_15__in1;
  wire [15:0] op_6_15__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_15(
    .in0(op_6_15__in0),
    .in1(op_6_15__in1),
    .out(op_6_15__out)
  );

  //Wire declarations for instance 'op_6_16' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_16__in0;
  wire [15:0] op_6_16__in1;
  wire [15:0] op_6_16__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_16(
    .in0(op_6_16__in0),
    .in1(op_6_16__in1),
    .out(op_6_16__out)
  );

  //Wire declarations for instance 'op_6_17' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_17__in0;
  wire [15:0] op_6_17__in1;
  wire [15:0] op_6_17__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_17(
    .in0(op_6_17__in0),
    .in1(op_6_17__in1),
    .out(op_6_17__out)
  );

  //Wire declarations for instance 'op_6_18' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_18__in0;
  wire [15:0] op_6_18__in1;
  wire [15:0] op_6_18__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_18(
    .in0(op_6_18__in0),
    .in1(op_6_18__in1),
    .out(op_6_18__out)
  );

  //Wire declarations for instance 'op_6_19' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_19__in0;
  wire [15:0] op_6_19__in1;
  wire [15:0] op_6_19__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_19(
    .in0(op_6_19__in0),
    .in1(op_6_19__in1),
    .out(op_6_19__out)
  );

  //Wire declarations for instance 'op_6_2' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_2__in0;
  wire [15:0] op_6_2__in1;
  wire [15:0] op_6_2__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_2(
    .in0(op_6_2__in0),
    .in1(op_6_2__in1),
    .out(op_6_2__out)
  );

  //Wire declarations for instance 'op_6_20' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_20__in0;
  wire [15:0] op_6_20__in1;
  wire [15:0] op_6_20__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_20(
    .in0(op_6_20__in0),
    .in1(op_6_20__in1),
    .out(op_6_20__out)
  );

  //Wire declarations for instance 'op_6_21' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_21__in0;
  wire [15:0] op_6_21__in1;
  wire [15:0] op_6_21__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_21(
    .in0(op_6_21__in0),
    .in1(op_6_21__in1),
    .out(op_6_21__out)
  );

  //Wire declarations for instance 'op_6_22' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_22__in0;
  wire [15:0] op_6_22__in1;
  wire [15:0] op_6_22__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_22(
    .in0(op_6_22__in0),
    .in1(op_6_22__in1),
    .out(op_6_22__out)
  );

  //Wire declarations for instance 'op_6_23' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_23__in0;
  wire [15:0] op_6_23__in1;
  wire [15:0] op_6_23__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_23(
    .in0(op_6_23__in0),
    .in1(op_6_23__in1),
    .out(op_6_23__out)
  );

  //Wire declarations for instance 'op_6_24' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_24__in0;
  wire [15:0] op_6_24__in1;
  wire [15:0] op_6_24__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_24(
    .in0(op_6_24__in0),
    .in1(op_6_24__in1),
    .out(op_6_24__out)
  );

  //Wire declarations for instance 'op_6_25' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_25__in0;
  wire [15:0] op_6_25__in1;
  wire [15:0] op_6_25__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_25(
    .in0(op_6_25__in0),
    .in1(op_6_25__in1),
    .out(op_6_25__out)
  );

  //Wire declarations for instance 'op_6_26' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_26__in0;
  wire [15:0] op_6_26__in1;
  wire [15:0] op_6_26__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_26(
    .in0(op_6_26__in0),
    .in1(op_6_26__in1),
    .out(op_6_26__out)
  );

  //Wire declarations for instance 'op_6_27' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_27__in0;
  wire [15:0] op_6_27__in1;
  wire [15:0] op_6_27__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_27(
    .in0(op_6_27__in0),
    .in1(op_6_27__in1),
    .out(op_6_27__out)
  );

  //Wire declarations for instance 'op_6_28' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_28__in0;
  wire [15:0] op_6_28__in1;
  wire [15:0] op_6_28__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_28(
    .in0(op_6_28__in0),
    .in1(op_6_28__in1),
    .out(op_6_28__out)
  );

  //Wire declarations for instance 'op_6_29' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_29__in0;
  wire [15:0] op_6_29__in1;
  wire [15:0] op_6_29__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_29(
    .in0(op_6_29__in0),
    .in1(op_6_29__in1),
    .out(op_6_29__out)
  );

  //Wire declarations for instance 'op_6_3' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_3__in0;
  wire [15:0] op_6_3__in1;
  wire [15:0] op_6_3__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_3(
    .in0(op_6_3__in0),
    .in1(op_6_3__in1),
    .out(op_6_3__out)
  );

  //Wire declarations for instance 'op_6_30' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_30__in0;
  wire [15:0] op_6_30__in1;
  wire [15:0] op_6_30__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_30(
    .in0(op_6_30__in0),
    .in1(op_6_30__in1),
    .out(op_6_30__out)
  );

  //Wire declarations for instance 'op_6_31' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_31__in0;
  wire [15:0] op_6_31__in1;
  wire [15:0] op_6_31__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_31(
    .in0(op_6_31__in0),
    .in1(op_6_31__in1),
    .out(op_6_31__out)
  );

  //Wire declarations for instance 'op_6_32' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_32__in0;
  wire [15:0] op_6_32__in1;
  wire [15:0] op_6_32__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_32(
    .in0(op_6_32__in0),
    .in1(op_6_32__in1),
    .out(op_6_32__out)
  );

  //Wire declarations for instance 'op_6_33' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_33__in0;
  wire [15:0] op_6_33__in1;
  wire [15:0] op_6_33__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_33(
    .in0(op_6_33__in0),
    .in1(op_6_33__in1),
    .out(op_6_33__out)
  );

  //Wire declarations for instance 'op_6_34' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_34__in0;
  wire [15:0] op_6_34__in1;
  wire [15:0] op_6_34__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_34(
    .in0(op_6_34__in0),
    .in1(op_6_34__in1),
    .out(op_6_34__out)
  );

  //Wire declarations for instance 'op_6_35' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_35__in0;
  wire [15:0] op_6_35__in1;
  wire [15:0] op_6_35__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_35(
    .in0(op_6_35__in0),
    .in1(op_6_35__in1),
    .out(op_6_35__out)
  );

  //Wire declarations for instance 'op_6_36' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_36__in0;
  wire [15:0] op_6_36__in1;
  wire [15:0] op_6_36__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_36(
    .in0(op_6_36__in0),
    .in1(op_6_36__in1),
    .out(op_6_36__out)
  );

  //Wire declarations for instance 'op_6_37' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_37__in0;
  wire [15:0] op_6_37__in1;
  wire [15:0] op_6_37__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_37(
    .in0(op_6_37__in0),
    .in1(op_6_37__in1),
    .out(op_6_37__out)
  );

  //Wire declarations for instance 'op_6_38' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_38__in0;
  wire [15:0] op_6_38__in1;
  wire [15:0] op_6_38__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_38(
    .in0(op_6_38__in0),
    .in1(op_6_38__in1),
    .out(op_6_38__out)
  );

  //Wire declarations for instance 'op_6_39' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_39__in0;
  wire [15:0] op_6_39__in1;
  wire [15:0] op_6_39__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_39(
    .in0(op_6_39__in0),
    .in1(op_6_39__in1),
    .out(op_6_39__out)
  );

  //Wire declarations for instance 'op_6_4' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_4__in0;
  wire [15:0] op_6_4__in1;
  wire [15:0] op_6_4__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_4(
    .in0(op_6_4__in0),
    .in1(op_6_4__in1),
    .out(op_6_4__out)
  );

  //Wire declarations for instance 'op_6_40' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_40__in0;
  wire [15:0] op_6_40__in1;
  wire [15:0] op_6_40__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_40(
    .in0(op_6_40__in0),
    .in1(op_6_40__in1),
    .out(op_6_40__out)
  );

  //Wire declarations for instance 'op_6_41' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_41__in0;
  wire [15:0] op_6_41__in1;
  wire [15:0] op_6_41__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_41(
    .in0(op_6_41__in0),
    .in1(op_6_41__in1),
    .out(op_6_41__out)
  );

  //Wire declarations for instance 'op_6_42' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_42__in0;
  wire [15:0] op_6_42__in1;
  wire [15:0] op_6_42__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_42(
    .in0(op_6_42__in0),
    .in1(op_6_42__in1),
    .out(op_6_42__out)
  );

  //Wire declarations for instance 'op_6_43' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_43__in0;
  wire [15:0] op_6_43__in1;
  wire [15:0] op_6_43__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_43(
    .in0(op_6_43__in0),
    .in1(op_6_43__in1),
    .out(op_6_43__out)
  );

  //Wire declarations for instance 'op_6_44' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_44__in0;
  wire [15:0] op_6_44__in1;
  wire [15:0] op_6_44__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_44(
    .in0(op_6_44__in0),
    .in1(op_6_44__in1),
    .out(op_6_44__out)
  );

  //Wire declarations for instance 'op_6_45' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_45__in0;
  wire [15:0] op_6_45__in1;
  wire [15:0] op_6_45__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_45(
    .in0(op_6_45__in0),
    .in1(op_6_45__in1),
    .out(op_6_45__out)
  );

  //Wire declarations for instance 'op_6_46' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_46__in0;
  wire [15:0] op_6_46__in1;
  wire [15:0] op_6_46__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_46(
    .in0(op_6_46__in0),
    .in1(op_6_46__in1),
    .out(op_6_46__out)
  );

  //Wire declarations for instance 'op_6_47' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_47__in0;
  wire [15:0] op_6_47__in1;
  wire [15:0] op_6_47__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_47(
    .in0(op_6_47__in0),
    .in1(op_6_47__in1),
    .out(op_6_47__out)
  );

  //Wire declarations for instance 'op_6_48' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_48__in0;
  wire [15:0] op_6_48__in1;
  wire [15:0] op_6_48__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_48(
    .in0(op_6_48__in0),
    .in1(op_6_48__in1),
    .out(op_6_48__out)
  );

  //Wire declarations for instance 'op_6_49' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_49__in0;
  wire [15:0] op_6_49__in1;
  wire [15:0] op_6_49__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_49(
    .in0(op_6_49__in0),
    .in1(op_6_49__in1),
    .out(op_6_49__out)
  );

  //Wire declarations for instance 'op_6_5' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_5__in0;
  wire [15:0] op_6_5__in1;
  wire [15:0] op_6_5__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_5(
    .in0(op_6_5__in0),
    .in1(op_6_5__in1),
    .out(op_6_5__out)
  );

  //Wire declarations for instance 'op_6_50' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_50__in0;
  wire [15:0] op_6_50__in1;
  wire [15:0] op_6_50__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_50(
    .in0(op_6_50__in0),
    .in1(op_6_50__in1),
    .out(op_6_50__out)
  );

  //Wire declarations for instance 'op_6_51' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_51__in0;
  wire [15:0] op_6_51__in1;
  wire [15:0] op_6_51__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_51(
    .in0(op_6_51__in0),
    .in1(op_6_51__in1),
    .out(op_6_51__out)
  );

  //Wire declarations for instance 'op_6_52' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_52__in0;
  wire [15:0] op_6_52__in1;
  wire [15:0] op_6_52__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_52(
    .in0(op_6_52__in0),
    .in1(op_6_52__in1),
    .out(op_6_52__out)
  );

  //Wire declarations for instance 'op_6_53' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_53__in0;
  wire [15:0] op_6_53__in1;
  wire [15:0] op_6_53__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_53(
    .in0(op_6_53__in0),
    .in1(op_6_53__in1),
    .out(op_6_53__out)
  );

  //Wire declarations for instance 'op_6_54' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_54__in0;
  wire [15:0] op_6_54__in1;
  wire [15:0] op_6_54__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_54(
    .in0(op_6_54__in0),
    .in1(op_6_54__in1),
    .out(op_6_54__out)
  );

  //Wire declarations for instance 'op_6_55' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_55__in0;
  wire [15:0] op_6_55__in1;
  wire [15:0] op_6_55__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_55(
    .in0(op_6_55__in0),
    .in1(op_6_55__in1),
    .out(op_6_55__out)
  );

  //Wire declarations for instance 'op_6_56' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_56__in0;
  wire [15:0] op_6_56__in1;
  wire [15:0] op_6_56__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_56(
    .in0(op_6_56__in0),
    .in1(op_6_56__in1),
    .out(op_6_56__out)
  );

  //Wire declarations for instance 'op_6_57' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_57__in0;
  wire [15:0] op_6_57__in1;
  wire [15:0] op_6_57__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_57(
    .in0(op_6_57__in0),
    .in1(op_6_57__in1),
    .out(op_6_57__out)
  );

  //Wire declarations for instance 'op_6_58' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_58__in0;
  wire [15:0] op_6_58__in1;
  wire [15:0] op_6_58__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_58(
    .in0(op_6_58__in0),
    .in1(op_6_58__in1),
    .out(op_6_58__out)
  );

  //Wire declarations for instance 'op_6_59' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_59__in0;
  wire [15:0] op_6_59__in1;
  wire [15:0] op_6_59__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_59(
    .in0(op_6_59__in0),
    .in1(op_6_59__in1),
    .out(op_6_59__out)
  );

  //Wire declarations for instance 'op_6_6' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_6__in0;
  wire [15:0] op_6_6__in1;
  wire [15:0] op_6_6__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_6(
    .in0(op_6_6__in0),
    .in1(op_6_6__in1),
    .out(op_6_6__out)
  );

  //Wire declarations for instance 'op_6_60' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_60__in0;
  wire [15:0] op_6_60__in1;
  wire [15:0] op_6_60__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_60(
    .in0(op_6_60__in0),
    .in1(op_6_60__in1),
    .out(op_6_60__out)
  );

  //Wire declarations for instance 'op_6_61' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_61__in0;
  wire [15:0] op_6_61__in1;
  wire [15:0] op_6_61__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_61(
    .in0(op_6_61__in0),
    .in1(op_6_61__in1),
    .out(op_6_61__out)
  );

  //Wire declarations for instance 'op_6_62' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_62__in0;
  wire [15:0] op_6_62__in1;
  wire [15:0] op_6_62__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_62(
    .in0(op_6_62__in0),
    .in1(op_6_62__in1),
    .out(op_6_62__out)
  );

  //Wire declarations for instance 'op_6_63' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_63__in0;
  wire [15:0] op_6_63__in1;
  wire [15:0] op_6_63__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_63(
    .in0(op_6_63__in0),
    .in1(op_6_63__in1),
    .out(op_6_63__out)
  );

  //Wire declarations for instance 'op_6_7' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_7__in0;
  wire [15:0] op_6_7__in1;
  wire [15:0] op_6_7__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_7(
    .in0(op_6_7__in0),
    .in1(op_6_7__in1),
    .out(op_6_7__out)
  );

  //Wire declarations for instance 'op_6_8' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_8__in0;
  wire [15:0] op_6_8__in1;
  wire [15:0] op_6_8__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_8(
    .in0(op_6_8__in0),
    .in1(op_6_8__in1),
    .out(op_6_8__out)
  );

  //Wire declarations for instance 'op_6_9' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_6_9__in0;
  wire [15:0] op_6_9__in1;
  wire [15:0] op_6_9__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_6_9(
    .in0(op_6_9__in0),
    .in1(op_6_9__in1),
    .out(op_6_9__out)
  );

  //Wire declarations for instance 'op_7_0' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_0__in0;
  wire [15:0] op_7_0__in1;
  wire [15:0] op_7_0__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_0(
    .in0(op_7_0__in0),
    .in1(op_7_0__in1),
    .out(op_7_0__out)
  );

  //Wire declarations for instance 'op_7_1' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_1__in0;
  wire [15:0] op_7_1__in1;
  wire [15:0] op_7_1__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_1(
    .in0(op_7_1__in0),
    .in1(op_7_1__in1),
    .out(op_7_1__out)
  );

  //Wire declarations for instance 'op_7_10' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_10__in0;
  wire [15:0] op_7_10__in1;
  wire [15:0] op_7_10__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_10(
    .in0(op_7_10__in0),
    .in1(op_7_10__in1),
    .out(op_7_10__out)
  );

  //Wire declarations for instance 'op_7_100' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_100__in0;
  wire [15:0] op_7_100__in1;
  wire [15:0] op_7_100__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_100(
    .in0(op_7_100__in0),
    .in1(op_7_100__in1),
    .out(op_7_100__out)
  );

  //Wire declarations for instance 'op_7_101' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_101__in0;
  wire [15:0] op_7_101__in1;
  wire [15:0] op_7_101__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_101(
    .in0(op_7_101__in0),
    .in1(op_7_101__in1),
    .out(op_7_101__out)
  );

  //Wire declarations for instance 'op_7_102' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_102__in0;
  wire [15:0] op_7_102__in1;
  wire [15:0] op_7_102__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_102(
    .in0(op_7_102__in0),
    .in1(op_7_102__in1),
    .out(op_7_102__out)
  );

  //Wire declarations for instance 'op_7_103' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_103__in0;
  wire [15:0] op_7_103__in1;
  wire [15:0] op_7_103__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_103(
    .in0(op_7_103__in0),
    .in1(op_7_103__in1),
    .out(op_7_103__out)
  );

  //Wire declarations for instance 'op_7_104' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_104__in0;
  wire [15:0] op_7_104__in1;
  wire [15:0] op_7_104__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_104(
    .in0(op_7_104__in0),
    .in1(op_7_104__in1),
    .out(op_7_104__out)
  );

  //Wire declarations for instance 'op_7_105' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_105__in0;
  wire [15:0] op_7_105__in1;
  wire [15:0] op_7_105__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_105(
    .in0(op_7_105__in0),
    .in1(op_7_105__in1),
    .out(op_7_105__out)
  );

  //Wire declarations for instance 'op_7_106' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_106__in0;
  wire [15:0] op_7_106__in1;
  wire [15:0] op_7_106__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_106(
    .in0(op_7_106__in0),
    .in1(op_7_106__in1),
    .out(op_7_106__out)
  );

  //Wire declarations for instance 'op_7_107' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_107__in0;
  wire [15:0] op_7_107__in1;
  wire [15:0] op_7_107__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_107(
    .in0(op_7_107__in0),
    .in1(op_7_107__in1),
    .out(op_7_107__out)
  );

  //Wire declarations for instance 'op_7_108' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_108__in0;
  wire [15:0] op_7_108__in1;
  wire [15:0] op_7_108__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_108(
    .in0(op_7_108__in0),
    .in1(op_7_108__in1),
    .out(op_7_108__out)
  );

  //Wire declarations for instance 'op_7_109' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_109__in0;
  wire [15:0] op_7_109__in1;
  wire [15:0] op_7_109__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_109(
    .in0(op_7_109__in0),
    .in1(op_7_109__in1),
    .out(op_7_109__out)
  );

  //Wire declarations for instance 'op_7_11' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_11__in0;
  wire [15:0] op_7_11__in1;
  wire [15:0] op_7_11__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_11(
    .in0(op_7_11__in0),
    .in1(op_7_11__in1),
    .out(op_7_11__out)
  );

  //Wire declarations for instance 'op_7_110' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_110__in0;
  wire [15:0] op_7_110__in1;
  wire [15:0] op_7_110__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_110(
    .in0(op_7_110__in0),
    .in1(op_7_110__in1),
    .out(op_7_110__out)
  );

  //Wire declarations for instance 'op_7_111' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_111__in0;
  wire [15:0] op_7_111__in1;
  wire [15:0] op_7_111__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_111(
    .in0(op_7_111__in0),
    .in1(op_7_111__in1),
    .out(op_7_111__out)
  );

  //Wire declarations for instance 'op_7_112' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_112__in0;
  wire [15:0] op_7_112__in1;
  wire [15:0] op_7_112__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_112(
    .in0(op_7_112__in0),
    .in1(op_7_112__in1),
    .out(op_7_112__out)
  );

  //Wire declarations for instance 'op_7_113' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_113__in0;
  wire [15:0] op_7_113__in1;
  wire [15:0] op_7_113__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_113(
    .in0(op_7_113__in0),
    .in1(op_7_113__in1),
    .out(op_7_113__out)
  );

  //Wire declarations for instance 'op_7_114' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_114__in0;
  wire [15:0] op_7_114__in1;
  wire [15:0] op_7_114__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_114(
    .in0(op_7_114__in0),
    .in1(op_7_114__in1),
    .out(op_7_114__out)
  );

  //Wire declarations for instance 'op_7_115' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_115__in0;
  wire [15:0] op_7_115__in1;
  wire [15:0] op_7_115__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_115(
    .in0(op_7_115__in0),
    .in1(op_7_115__in1),
    .out(op_7_115__out)
  );

  //Wire declarations for instance 'op_7_116' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_116__in0;
  wire [15:0] op_7_116__in1;
  wire [15:0] op_7_116__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_116(
    .in0(op_7_116__in0),
    .in1(op_7_116__in1),
    .out(op_7_116__out)
  );

  //Wire declarations for instance 'op_7_117' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_117__in0;
  wire [15:0] op_7_117__in1;
  wire [15:0] op_7_117__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_117(
    .in0(op_7_117__in0),
    .in1(op_7_117__in1),
    .out(op_7_117__out)
  );

  //Wire declarations for instance 'op_7_118' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_118__in0;
  wire [15:0] op_7_118__in1;
  wire [15:0] op_7_118__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_118(
    .in0(op_7_118__in0),
    .in1(op_7_118__in1),
    .out(op_7_118__out)
  );

  //Wire declarations for instance 'op_7_119' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_119__in0;
  wire [15:0] op_7_119__in1;
  wire [15:0] op_7_119__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_119(
    .in0(op_7_119__in0),
    .in1(op_7_119__in1),
    .out(op_7_119__out)
  );

  //Wire declarations for instance 'op_7_12' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_12__in0;
  wire [15:0] op_7_12__in1;
  wire [15:0] op_7_12__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_12(
    .in0(op_7_12__in0),
    .in1(op_7_12__in1),
    .out(op_7_12__out)
  );

  //Wire declarations for instance 'op_7_120' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_120__in0;
  wire [15:0] op_7_120__in1;
  wire [15:0] op_7_120__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_120(
    .in0(op_7_120__in0),
    .in1(op_7_120__in1),
    .out(op_7_120__out)
  );

  //Wire declarations for instance 'op_7_121' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_121__in0;
  wire [15:0] op_7_121__in1;
  wire [15:0] op_7_121__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_121(
    .in0(op_7_121__in0),
    .in1(op_7_121__in1),
    .out(op_7_121__out)
  );

  //Wire declarations for instance 'op_7_122' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_122__in0;
  wire [15:0] op_7_122__in1;
  wire [15:0] op_7_122__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_122(
    .in0(op_7_122__in0),
    .in1(op_7_122__in1),
    .out(op_7_122__out)
  );

  //Wire declarations for instance 'op_7_123' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_123__in0;
  wire [15:0] op_7_123__in1;
  wire [15:0] op_7_123__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_123(
    .in0(op_7_123__in0),
    .in1(op_7_123__in1),
    .out(op_7_123__out)
  );

  //Wire declarations for instance 'op_7_124' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_124__in0;
  wire [15:0] op_7_124__in1;
  wire [15:0] op_7_124__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_124(
    .in0(op_7_124__in0),
    .in1(op_7_124__in1),
    .out(op_7_124__out)
  );

  //Wire declarations for instance 'op_7_125' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_125__in0;
  wire [15:0] op_7_125__in1;
  wire [15:0] op_7_125__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_125(
    .in0(op_7_125__in0),
    .in1(op_7_125__in1),
    .out(op_7_125__out)
  );

  //Wire declarations for instance 'op_7_126' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_126__in0;
  wire [15:0] op_7_126__in1;
  wire [15:0] op_7_126__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_126(
    .in0(op_7_126__in0),
    .in1(op_7_126__in1),
    .out(op_7_126__out)
  );

  //Wire declarations for instance 'op_7_127' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_127__in0;
  wire [15:0] op_7_127__in1;
  wire [15:0] op_7_127__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_127(
    .in0(op_7_127__in0),
    .in1(op_7_127__in1),
    .out(op_7_127__out)
  );

  //Wire declarations for instance 'op_7_13' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_13__in0;
  wire [15:0] op_7_13__in1;
  wire [15:0] op_7_13__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_13(
    .in0(op_7_13__in0),
    .in1(op_7_13__in1),
    .out(op_7_13__out)
  );

  //Wire declarations for instance 'op_7_14' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_14__in0;
  wire [15:0] op_7_14__in1;
  wire [15:0] op_7_14__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_14(
    .in0(op_7_14__in0),
    .in1(op_7_14__in1),
    .out(op_7_14__out)
  );

  //Wire declarations for instance 'op_7_15' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_15__in0;
  wire [15:0] op_7_15__in1;
  wire [15:0] op_7_15__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_15(
    .in0(op_7_15__in0),
    .in1(op_7_15__in1),
    .out(op_7_15__out)
  );

  //Wire declarations for instance 'op_7_16' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_16__in0;
  wire [15:0] op_7_16__in1;
  wire [15:0] op_7_16__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_16(
    .in0(op_7_16__in0),
    .in1(op_7_16__in1),
    .out(op_7_16__out)
  );

  //Wire declarations for instance 'op_7_17' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_17__in0;
  wire [15:0] op_7_17__in1;
  wire [15:0] op_7_17__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_17(
    .in0(op_7_17__in0),
    .in1(op_7_17__in1),
    .out(op_7_17__out)
  );

  //Wire declarations for instance 'op_7_18' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_18__in0;
  wire [15:0] op_7_18__in1;
  wire [15:0] op_7_18__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_18(
    .in0(op_7_18__in0),
    .in1(op_7_18__in1),
    .out(op_7_18__out)
  );

  //Wire declarations for instance 'op_7_19' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_19__in0;
  wire [15:0] op_7_19__in1;
  wire [15:0] op_7_19__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_19(
    .in0(op_7_19__in0),
    .in1(op_7_19__in1),
    .out(op_7_19__out)
  );

  //Wire declarations for instance 'op_7_2' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_2__in0;
  wire [15:0] op_7_2__in1;
  wire [15:0] op_7_2__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_2(
    .in0(op_7_2__in0),
    .in1(op_7_2__in1),
    .out(op_7_2__out)
  );

  //Wire declarations for instance 'op_7_20' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_20__in0;
  wire [15:0] op_7_20__in1;
  wire [15:0] op_7_20__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_20(
    .in0(op_7_20__in0),
    .in1(op_7_20__in1),
    .out(op_7_20__out)
  );

  //Wire declarations for instance 'op_7_21' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_21__in0;
  wire [15:0] op_7_21__in1;
  wire [15:0] op_7_21__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_21(
    .in0(op_7_21__in0),
    .in1(op_7_21__in1),
    .out(op_7_21__out)
  );

  //Wire declarations for instance 'op_7_22' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_22__in0;
  wire [15:0] op_7_22__in1;
  wire [15:0] op_7_22__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_22(
    .in0(op_7_22__in0),
    .in1(op_7_22__in1),
    .out(op_7_22__out)
  );

  //Wire declarations for instance 'op_7_23' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_23__in0;
  wire [15:0] op_7_23__in1;
  wire [15:0] op_7_23__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_23(
    .in0(op_7_23__in0),
    .in1(op_7_23__in1),
    .out(op_7_23__out)
  );

  //Wire declarations for instance 'op_7_24' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_24__in0;
  wire [15:0] op_7_24__in1;
  wire [15:0] op_7_24__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_24(
    .in0(op_7_24__in0),
    .in1(op_7_24__in1),
    .out(op_7_24__out)
  );

  //Wire declarations for instance 'op_7_25' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_25__in0;
  wire [15:0] op_7_25__in1;
  wire [15:0] op_7_25__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_25(
    .in0(op_7_25__in0),
    .in1(op_7_25__in1),
    .out(op_7_25__out)
  );

  //Wire declarations for instance 'op_7_26' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_26__in0;
  wire [15:0] op_7_26__in1;
  wire [15:0] op_7_26__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_26(
    .in0(op_7_26__in0),
    .in1(op_7_26__in1),
    .out(op_7_26__out)
  );

  //Wire declarations for instance 'op_7_27' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_27__in0;
  wire [15:0] op_7_27__in1;
  wire [15:0] op_7_27__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_27(
    .in0(op_7_27__in0),
    .in1(op_7_27__in1),
    .out(op_7_27__out)
  );

  //Wire declarations for instance 'op_7_28' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_28__in0;
  wire [15:0] op_7_28__in1;
  wire [15:0] op_7_28__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_28(
    .in0(op_7_28__in0),
    .in1(op_7_28__in1),
    .out(op_7_28__out)
  );

  //Wire declarations for instance 'op_7_29' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_29__in0;
  wire [15:0] op_7_29__in1;
  wire [15:0] op_7_29__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_29(
    .in0(op_7_29__in0),
    .in1(op_7_29__in1),
    .out(op_7_29__out)
  );

  //Wire declarations for instance 'op_7_3' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_3__in0;
  wire [15:0] op_7_3__in1;
  wire [15:0] op_7_3__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_3(
    .in0(op_7_3__in0),
    .in1(op_7_3__in1),
    .out(op_7_3__out)
  );

  //Wire declarations for instance 'op_7_30' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_30__in0;
  wire [15:0] op_7_30__in1;
  wire [15:0] op_7_30__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_30(
    .in0(op_7_30__in0),
    .in1(op_7_30__in1),
    .out(op_7_30__out)
  );

  //Wire declarations for instance 'op_7_31' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_31__in0;
  wire [15:0] op_7_31__in1;
  wire [15:0] op_7_31__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_31(
    .in0(op_7_31__in0),
    .in1(op_7_31__in1),
    .out(op_7_31__out)
  );

  //Wire declarations for instance 'op_7_32' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_32__in0;
  wire [15:0] op_7_32__in1;
  wire [15:0] op_7_32__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_32(
    .in0(op_7_32__in0),
    .in1(op_7_32__in1),
    .out(op_7_32__out)
  );

  //Wire declarations for instance 'op_7_33' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_33__in0;
  wire [15:0] op_7_33__in1;
  wire [15:0] op_7_33__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_33(
    .in0(op_7_33__in0),
    .in1(op_7_33__in1),
    .out(op_7_33__out)
  );

  //Wire declarations for instance 'op_7_34' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_34__in0;
  wire [15:0] op_7_34__in1;
  wire [15:0] op_7_34__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_34(
    .in0(op_7_34__in0),
    .in1(op_7_34__in1),
    .out(op_7_34__out)
  );

  //Wire declarations for instance 'op_7_35' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_35__in0;
  wire [15:0] op_7_35__in1;
  wire [15:0] op_7_35__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_35(
    .in0(op_7_35__in0),
    .in1(op_7_35__in1),
    .out(op_7_35__out)
  );

  //Wire declarations for instance 'op_7_36' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_36__in0;
  wire [15:0] op_7_36__in1;
  wire [15:0] op_7_36__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_36(
    .in0(op_7_36__in0),
    .in1(op_7_36__in1),
    .out(op_7_36__out)
  );

  //Wire declarations for instance 'op_7_37' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_37__in0;
  wire [15:0] op_7_37__in1;
  wire [15:0] op_7_37__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_37(
    .in0(op_7_37__in0),
    .in1(op_7_37__in1),
    .out(op_7_37__out)
  );

  //Wire declarations for instance 'op_7_38' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_38__in0;
  wire [15:0] op_7_38__in1;
  wire [15:0] op_7_38__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_38(
    .in0(op_7_38__in0),
    .in1(op_7_38__in1),
    .out(op_7_38__out)
  );

  //Wire declarations for instance 'op_7_39' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_39__in0;
  wire [15:0] op_7_39__in1;
  wire [15:0] op_7_39__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_39(
    .in0(op_7_39__in0),
    .in1(op_7_39__in1),
    .out(op_7_39__out)
  );

  //Wire declarations for instance 'op_7_4' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_4__in0;
  wire [15:0] op_7_4__in1;
  wire [15:0] op_7_4__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_4(
    .in0(op_7_4__in0),
    .in1(op_7_4__in1),
    .out(op_7_4__out)
  );

  //Wire declarations for instance 'op_7_40' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_40__in0;
  wire [15:0] op_7_40__in1;
  wire [15:0] op_7_40__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_40(
    .in0(op_7_40__in0),
    .in1(op_7_40__in1),
    .out(op_7_40__out)
  );

  //Wire declarations for instance 'op_7_41' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_41__in0;
  wire [15:0] op_7_41__in1;
  wire [15:0] op_7_41__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_41(
    .in0(op_7_41__in0),
    .in1(op_7_41__in1),
    .out(op_7_41__out)
  );

  //Wire declarations for instance 'op_7_42' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_42__in0;
  wire [15:0] op_7_42__in1;
  wire [15:0] op_7_42__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_42(
    .in0(op_7_42__in0),
    .in1(op_7_42__in1),
    .out(op_7_42__out)
  );

  //Wire declarations for instance 'op_7_43' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_43__in0;
  wire [15:0] op_7_43__in1;
  wire [15:0] op_7_43__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_43(
    .in0(op_7_43__in0),
    .in1(op_7_43__in1),
    .out(op_7_43__out)
  );

  //Wire declarations for instance 'op_7_44' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_44__in0;
  wire [15:0] op_7_44__in1;
  wire [15:0] op_7_44__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_44(
    .in0(op_7_44__in0),
    .in1(op_7_44__in1),
    .out(op_7_44__out)
  );

  //Wire declarations for instance 'op_7_45' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_45__in0;
  wire [15:0] op_7_45__in1;
  wire [15:0] op_7_45__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_45(
    .in0(op_7_45__in0),
    .in1(op_7_45__in1),
    .out(op_7_45__out)
  );

  //Wire declarations for instance 'op_7_46' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_46__in0;
  wire [15:0] op_7_46__in1;
  wire [15:0] op_7_46__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_46(
    .in0(op_7_46__in0),
    .in1(op_7_46__in1),
    .out(op_7_46__out)
  );

  //Wire declarations for instance 'op_7_47' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_47__in0;
  wire [15:0] op_7_47__in1;
  wire [15:0] op_7_47__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_47(
    .in0(op_7_47__in0),
    .in1(op_7_47__in1),
    .out(op_7_47__out)
  );

  //Wire declarations for instance 'op_7_48' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_48__in0;
  wire [15:0] op_7_48__in1;
  wire [15:0] op_7_48__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_48(
    .in0(op_7_48__in0),
    .in1(op_7_48__in1),
    .out(op_7_48__out)
  );

  //Wire declarations for instance 'op_7_49' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_49__in0;
  wire [15:0] op_7_49__in1;
  wire [15:0] op_7_49__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_49(
    .in0(op_7_49__in0),
    .in1(op_7_49__in1),
    .out(op_7_49__out)
  );

  //Wire declarations for instance 'op_7_5' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_5__in0;
  wire [15:0] op_7_5__in1;
  wire [15:0] op_7_5__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_5(
    .in0(op_7_5__in0),
    .in1(op_7_5__in1),
    .out(op_7_5__out)
  );

  //Wire declarations for instance 'op_7_50' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_50__in0;
  wire [15:0] op_7_50__in1;
  wire [15:0] op_7_50__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_50(
    .in0(op_7_50__in0),
    .in1(op_7_50__in1),
    .out(op_7_50__out)
  );

  //Wire declarations for instance 'op_7_51' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_51__in0;
  wire [15:0] op_7_51__in1;
  wire [15:0] op_7_51__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_51(
    .in0(op_7_51__in0),
    .in1(op_7_51__in1),
    .out(op_7_51__out)
  );

  //Wire declarations for instance 'op_7_52' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_52__in0;
  wire [15:0] op_7_52__in1;
  wire [15:0] op_7_52__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_52(
    .in0(op_7_52__in0),
    .in1(op_7_52__in1),
    .out(op_7_52__out)
  );

  //Wire declarations for instance 'op_7_53' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_53__in0;
  wire [15:0] op_7_53__in1;
  wire [15:0] op_7_53__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_53(
    .in0(op_7_53__in0),
    .in1(op_7_53__in1),
    .out(op_7_53__out)
  );

  //Wire declarations for instance 'op_7_54' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_54__in0;
  wire [15:0] op_7_54__in1;
  wire [15:0] op_7_54__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_54(
    .in0(op_7_54__in0),
    .in1(op_7_54__in1),
    .out(op_7_54__out)
  );

  //Wire declarations for instance 'op_7_55' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_55__in0;
  wire [15:0] op_7_55__in1;
  wire [15:0] op_7_55__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_55(
    .in0(op_7_55__in0),
    .in1(op_7_55__in1),
    .out(op_7_55__out)
  );

  //Wire declarations for instance 'op_7_56' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_56__in0;
  wire [15:0] op_7_56__in1;
  wire [15:0] op_7_56__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_56(
    .in0(op_7_56__in0),
    .in1(op_7_56__in1),
    .out(op_7_56__out)
  );

  //Wire declarations for instance 'op_7_57' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_57__in0;
  wire [15:0] op_7_57__in1;
  wire [15:0] op_7_57__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_57(
    .in0(op_7_57__in0),
    .in1(op_7_57__in1),
    .out(op_7_57__out)
  );

  //Wire declarations for instance 'op_7_58' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_58__in0;
  wire [15:0] op_7_58__in1;
  wire [15:0] op_7_58__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_58(
    .in0(op_7_58__in0),
    .in1(op_7_58__in1),
    .out(op_7_58__out)
  );

  //Wire declarations for instance 'op_7_59' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_59__in0;
  wire [15:0] op_7_59__in1;
  wire [15:0] op_7_59__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_59(
    .in0(op_7_59__in0),
    .in1(op_7_59__in1),
    .out(op_7_59__out)
  );

  //Wire declarations for instance 'op_7_6' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_6__in0;
  wire [15:0] op_7_6__in1;
  wire [15:0] op_7_6__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_6(
    .in0(op_7_6__in0),
    .in1(op_7_6__in1),
    .out(op_7_6__out)
  );

  //Wire declarations for instance 'op_7_60' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_60__in0;
  wire [15:0] op_7_60__in1;
  wire [15:0] op_7_60__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_60(
    .in0(op_7_60__in0),
    .in1(op_7_60__in1),
    .out(op_7_60__out)
  );

  //Wire declarations for instance 'op_7_61' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_61__in0;
  wire [15:0] op_7_61__in1;
  wire [15:0] op_7_61__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_61(
    .in0(op_7_61__in0),
    .in1(op_7_61__in1),
    .out(op_7_61__out)
  );

  //Wire declarations for instance 'op_7_62' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_62__in0;
  wire [15:0] op_7_62__in1;
  wire [15:0] op_7_62__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_62(
    .in0(op_7_62__in0),
    .in1(op_7_62__in1),
    .out(op_7_62__out)
  );

  //Wire declarations for instance 'op_7_63' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_63__in0;
  wire [15:0] op_7_63__in1;
  wire [15:0] op_7_63__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_63(
    .in0(op_7_63__in0),
    .in1(op_7_63__in1),
    .out(op_7_63__out)
  );

  //Wire declarations for instance 'op_7_64' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_64__in0;
  wire [15:0] op_7_64__in1;
  wire [15:0] op_7_64__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_64(
    .in0(op_7_64__in0),
    .in1(op_7_64__in1),
    .out(op_7_64__out)
  );

  //Wire declarations for instance 'op_7_65' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_65__in0;
  wire [15:0] op_7_65__in1;
  wire [15:0] op_7_65__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_65(
    .in0(op_7_65__in0),
    .in1(op_7_65__in1),
    .out(op_7_65__out)
  );

  //Wire declarations for instance 'op_7_66' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_66__in0;
  wire [15:0] op_7_66__in1;
  wire [15:0] op_7_66__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_66(
    .in0(op_7_66__in0),
    .in1(op_7_66__in1),
    .out(op_7_66__out)
  );

  //Wire declarations for instance 'op_7_67' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_67__in0;
  wire [15:0] op_7_67__in1;
  wire [15:0] op_7_67__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_67(
    .in0(op_7_67__in0),
    .in1(op_7_67__in1),
    .out(op_7_67__out)
  );

  //Wire declarations for instance 'op_7_68' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_68__in0;
  wire [15:0] op_7_68__in1;
  wire [15:0] op_7_68__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_68(
    .in0(op_7_68__in0),
    .in1(op_7_68__in1),
    .out(op_7_68__out)
  );

  //Wire declarations for instance 'op_7_69' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_69__in0;
  wire [15:0] op_7_69__in1;
  wire [15:0] op_7_69__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_69(
    .in0(op_7_69__in0),
    .in1(op_7_69__in1),
    .out(op_7_69__out)
  );

  //Wire declarations for instance 'op_7_7' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_7__in0;
  wire [15:0] op_7_7__in1;
  wire [15:0] op_7_7__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_7(
    .in0(op_7_7__in0),
    .in1(op_7_7__in1),
    .out(op_7_7__out)
  );

  //Wire declarations for instance 'op_7_70' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_70__in0;
  wire [15:0] op_7_70__in1;
  wire [15:0] op_7_70__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_70(
    .in0(op_7_70__in0),
    .in1(op_7_70__in1),
    .out(op_7_70__out)
  );

  //Wire declarations for instance 'op_7_71' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_71__in0;
  wire [15:0] op_7_71__in1;
  wire [15:0] op_7_71__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_71(
    .in0(op_7_71__in0),
    .in1(op_7_71__in1),
    .out(op_7_71__out)
  );

  //Wire declarations for instance 'op_7_72' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_72__in0;
  wire [15:0] op_7_72__in1;
  wire [15:0] op_7_72__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_72(
    .in0(op_7_72__in0),
    .in1(op_7_72__in1),
    .out(op_7_72__out)
  );

  //Wire declarations for instance 'op_7_73' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_73__in0;
  wire [15:0] op_7_73__in1;
  wire [15:0] op_7_73__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_73(
    .in0(op_7_73__in0),
    .in1(op_7_73__in1),
    .out(op_7_73__out)
  );

  //Wire declarations for instance 'op_7_74' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_74__in0;
  wire [15:0] op_7_74__in1;
  wire [15:0] op_7_74__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_74(
    .in0(op_7_74__in0),
    .in1(op_7_74__in1),
    .out(op_7_74__out)
  );

  //Wire declarations for instance 'op_7_75' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_75__in0;
  wire [15:0] op_7_75__in1;
  wire [15:0] op_7_75__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_75(
    .in0(op_7_75__in0),
    .in1(op_7_75__in1),
    .out(op_7_75__out)
  );

  //Wire declarations for instance 'op_7_76' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_76__in0;
  wire [15:0] op_7_76__in1;
  wire [15:0] op_7_76__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_76(
    .in0(op_7_76__in0),
    .in1(op_7_76__in1),
    .out(op_7_76__out)
  );

  //Wire declarations for instance 'op_7_77' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_77__in0;
  wire [15:0] op_7_77__in1;
  wire [15:0] op_7_77__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_77(
    .in0(op_7_77__in0),
    .in1(op_7_77__in1),
    .out(op_7_77__out)
  );

  //Wire declarations for instance 'op_7_78' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_78__in0;
  wire [15:0] op_7_78__in1;
  wire [15:0] op_7_78__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_78(
    .in0(op_7_78__in0),
    .in1(op_7_78__in1),
    .out(op_7_78__out)
  );

  //Wire declarations for instance 'op_7_79' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_79__in0;
  wire [15:0] op_7_79__in1;
  wire [15:0] op_7_79__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_79(
    .in0(op_7_79__in0),
    .in1(op_7_79__in1),
    .out(op_7_79__out)
  );

  //Wire declarations for instance 'op_7_8' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_8__in0;
  wire [15:0] op_7_8__in1;
  wire [15:0] op_7_8__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_8(
    .in0(op_7_8__in0),
    .in1(op_7_8__in1),
    .out(op_7_8__out)
  );

  //Wire declarations for instance 'op_7_80' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_80__in0;
  wire [15:0] op_7_80__in1;
  wire [15:0] op_7_80__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_80(
    .in0(op_7_80__in0),
    .in1(op_7_80__in1),
    .out(op_7_80__out)
  );

  //Wire declarations for instance 'op_7_81' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_81__in0;
  wire [15:0] op_7_81__in1;
  wire [15:0] op_7_81__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_81(
    .in0(op_7_81__in0),
    .in1(op_7_81__in1),
    .out(op_7_81__out)
  );

  //Wire declarations for instance 'op_7_82' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_82__in0;
  wire [15:0] op_7_82__in1;
  wire [15:0] op_7_82__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_82(
    .in0(op_7_82__in0),
    .in1(op_7_82__in1),
    .out(op_7_82__out)
  );

  //Wire declarations for instance 'op_7_83' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_83__in0;
  wire [15:0] op_7_83__in1;
  wire [15:0] op_7_83__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_83(
    .in0(op_7_83__in0),
    .in1(op_7_83__in1),
    .out(op_7_83__out)
  );

  //Wire declarations for instance 'op_7_84' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_84__in0;
  wire [15:0] op_7_84__in1;
  wire [15:0] op_7_84__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_84(
    .in0(op_7_84__in0),
    .in1(op_7_84__in1),
    .out(op_7_84__out)
  );

  //Wire declarations for instance 'op_7_85' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_85__in0;
  wire [15:0] op_7_85__in1;
  wire [15:0] op_7_85__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_85(
    .in0(op_7_85__in0),
    .in1(op_7_85__in1),
    .out(op_7_85__out)
  );

  //Wire declarations for instance 'op_7_86' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_86__in0;
  wire [15:0] op_7_86__in1;
  wire [15:0] op_7_86__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_86(
    .in0(op_7_86__in0),
    .in1(op_7_86__in1),
    .out(op_7_86__out)
  );

  //Wire declarations for instance 'op_7_87' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_87__in0;
  wire [15:0] op_7_87__in1;
  wire [15:0] op_7_87__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_87(
    .in0(op_7_87__in0),
    .in1(op_7_87__in1),
    .out(op_7_87__out)
  );

  //Wire declarations for instance 'op_7_88' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_88__in0;
  wire [15:0] op_7_88__in1;
  wire [15:0] op_7_88__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_88(
    .in0(op_7_88__in0),
    .in1(op_7_88__in1),
    .out(op_7_88__out)
  );

  //Wire declarations for instance 'op_7_89' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_89__in0;
  wire [15:0] op_7_89__in1;
  wire [15:0] op_7_89__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_89(
    .in0(op_7_89__in0),
    .in1(op_7_89__in1),
    .out(op_7_89__out)
  );

  //Wire declarations for instance 'op_7_9' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_9__in0;
  wire [15:0] op_7_9__in1;
  wire [15:0] op_7_9__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_9(
    .in0(op_7_9__in0),
    .in1(op_7_9__in1),
    .out(op_7_9__out)
  );

  //Wire declarations for instance 'op_7_90' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_90__in0;
  wire [15:0] op_7_90__in1;
  wire [15:0] op_7_90__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_90(
    .in0(op_7_90__in0),
    .in1(op_7_90__in1),
    .out(op_7_90__out)
  );

  //Wire declarations for instance 'op_7_91' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_91__in0;
  wire [15:0] op_7_91__in1;
  wire [15:0] op_7_91__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_91(
    .in0(op_7_91__in0),
    .in1(op_7_91__in1),
    .out(op_7_91__out)
  );

  //Wire declarations for instance 'op_7_92' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_92__in0;
  wire [15:0] op_7_92__in1;
  wire [15:0] op_7_92__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_92(
    .in0(op_7_92__in0),
    .in1(op_7_92__in1),
    .out(op_7_92__out)
  );

  //Wire declarations for instance 'op_7_93' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_93__in0;
  wire [15:0] op_7_93__in1;
  wire [15:0] op_7_93__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_93(
    .in0(op_7_93__in0),
    .in1(op_7_93__in1),
    .out(op_7_93__out)
  );

  //Wire declarations for instance 'op_7_94' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_94__in0;
  wire [15:0] op_7_94__in1;
  wire [15:0] op_7_94__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_94(
    .in0(op_7_94__in0),
    .in1(op_7_94__in1),
    .out(op_7_94__out)
  );

  //Wire declarations for instance 'op_7_95' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_95__in0;
  wire [15:0] op_7_95__in1;
  wire [15:0] op_7_95__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_95(
    .in0(op_7_95__in0),
    .in1(op_7_95__in1),
    .out(op_7_95__out)
  );

  //Wire declarations for instance 'op_7_96' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_96__in0;
  wire [15:0] op_7_96__in1;
  wire [15:0] op_7_96__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_96(
    .in0(op_7_96__in0),
    .in1(op_7_96__in1),
    .out(op_7_96__out)
  );

  //Wire declarations for instance 'op_7_97' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_97__in0;
  wire [15:0] op_7_97__in1;
  wire [15:0] op_7_97__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_97(
    .in0(op_7_97__in0),
    .in1(op_7_97__in1),
    .out(op_7_97__out)
  );

  //Wire declarations for instance 'op_7_98' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_98__in0;
  wire [15:0] op_7_98__in1;
  wire [15:0] op_7_98__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_98(
    .in0(op_7_98__in0),
    .in1(op_7_98__in1),
    .out(op_7_98__out)
  );

  //Wire declarations for instance 'op_7_99' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_7_99__in0;
  wire [15:0] op_7_99__in1;
  wire [15:0] op_7_99__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_7_99(
    .in0(op_7_99__in0),
    .in1(op_7_99__in1),
    .out(op_7_99__out)
  );

  //Wire declarations for instance 'op_8_0' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_0__in0;
  wire [15:0] op_8_0__in1;
  wire [15:0] op_8_0__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_0(
    .in0(op_8_0__in0),
    .in1(op_8_0__in1),
    .out(op_8_0__out)
  );

  //Wire declarations for instance 'op_8_1' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_1__in0;
  wire [15:0] op_8_1__in1;
  wire [15:0] op_8_1__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_1(
    .in0(op_8_1__in0),
    .in1(op_8_1__in1),
    .out(op_8_1__out)
  );

  //Wire declarations for instance 'op_8_10' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_10__in0;
  wire [15:0] op_8_10__in1;
  wire [15:0] op_8_10__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_10(
    .in0(op_8_10__in0),
    .in1(op_8_10__in1),
    .out(op_8_10__out)
  );

  //Wire declarations for instance 'op_8_100' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_100__in0;
  wire [15:0] op_8_100__in1;
  wire [15:0] op_8_100__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_100(
    .in0(op_8_100__in0),
    .in1(op_8_100__in1),
    .out(op_8_100__out)
  );

  //Wire declarations for instance 'op_8_101' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_101__in0;
  wire [15:0] op_8_101__in1;
  wire [15:0] op_8_101__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_101(
    .in0(op_8_101__in0),
    .in1(op_8_101__in1),
    .out(op_8_101__out)
  );

  //Wire declarations for instance 'op_8_102' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_102__in0;
  wire [15:0] op_8_102__in1;
  wire [15:0] op_8_102__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_102(
    .in0(op_8_102__in0),
    .in1(op_8_102__in1),
    .out(op_8_102__out)
  );

  //Wire declarations for instance 'op_8_103' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_103__in0;
  wire [15:0] op_8_103__in1;
  wire [15:0] op_8_103__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_103(
    .in0(op_8_103__in0),
    .in1(op_8_103__in1),
    .out(op_8_103__out)
  );

  //Wire declarations for instance 'op_8_104' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_104__in0;
  wire [15:0] op_8_104__in1;
  wire [15:0] op_8_104__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_104(
    .in0(op_8_104__in0),
    .in1(op_8_104__in1),
    .out(op_8_104__out)
  );

  //Wire declarations for instance 'op_8_105' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_105__in0;
  wire [15:0] op_8_105__in1;
  wire [15:0] op_8_105__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_105(
    .in0(op_8_105__in0),
    .in1(op_8_105__in1),
    .out(op_8_105__out)
  );

  //Wire declarations for instance 'op_8_106' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_106__in0;
  wire [15:0] op_8_106__in1;
  wire [15:0] op_8_106__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_106(
    .in0(op_8_106__in0),
    .in1(op_8_106__in1),
    .out(op_8_106__out)
  );

  //Wire declarations for instance 'op_8_107' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_107__in0;
  wire [15:0] op_8_107__in1;
  wire [15:0] op_8_107__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_107(
    .in0(op_8_107__in0),
    .in1(op_8_107__in1),
    .out(op_8_107__out)
  );

  //Wire declarations for instance 'op_8_108' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_108__in0;
  wire [15:0] op_8_108__in1;
  wire [15:0] op_8_108__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_108(
    .in0(op_8_108__in0),
    .in1(op_8_108__in1),
    .out(op_8_108__out)
  );

  //Wire declarations for instance 'op_8_109' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_109__in0;
  wire [15:0] op_8_109__in1;
  wire [15:0] op_8_109__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_109(
    .in0(op_8_109__in0),
    .in1(op_8_109__in1),
    .out(op_8_109__out)
  );

  //Wire declarations for instance 'op_8_11' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_11__in0;
  wire [15:0] op_8_11__in1;
  wire [15:0] op_8_11__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_11(
    .in0(op_8_11__in0),
    .in1(op_8_11__in1),
    .out(op_8_11__out)
  );

  //Wire declarations for instance 'op_8_110' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_110__in0;
  wire [15:0] op_8_110__in1;
  wire [15:0] op_8_110__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_110(
    .in0(op_8_110__in0),
    .in1(op_8_110__in1),
    .out(op_8_110__out)
  );

  //Wire declarations for instance 'op_8_111' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_111__in0;
  wire [15:0] op_8_111__in1;
  wire [15:0] op_8_111__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_111(
    .in0(op_8_111__in0),
    .in1(op_8_111__in1),
    .out(op_8_111__out)
  );

  //Wire declarations for instance 'op_8_112' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_112__in0;
  wire [15:0] op_8_112__in1;
  wire [15:0] op_8_112__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_112(
    .in0(op_8_112__in0),
    .in1(op_8_112__in1),
    .out(op_8_112__out)
  );

  //Wire declarations for instance 'op_8_113' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_113__in0;
  wire [15:0] op_8_113__in1;
  wire [15:0] op_8_113__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_113(
    .in0(op_8_113__in0),
    .in1(op_8_113__in1),
    .out(op_8_113__out)
  );

  //Wire declarations for instance 'op_8_114' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_114__in0;
  wire [15:0] op_8_114__in1;
  wire [15:0] op_8_114__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_114(
    .in0(op_8_114__in0),
    .in1(op_8_114__in1),
    .out(op_8_114__out)
  );

  //Wire declarations for instance 'op_8_115' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_115__in0;
  wire [15:0] op_8_115__in1;
  wire [15:0] op_8_115__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_115(
    .in0(op_8_115__in0),
    .in1(op_8_115__in1),
    .out(op_8_115__out)
  );

  //Wire declarations for instance 'op_8_116' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_116__in0;
  wire [15:0] op_8_116__in1;
  wire [15:0] op_8_116__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_116(
    .in0(op_8_116__in0),
    .in1(op_8_116__in1),
    .out(op_8_116__out)
  );

  //Wire declarations for instance 'op_8_117' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_117__in0;
  wire [15:0] op_8_117__in1;
  wire [15:0] op_8_117__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_117(
    .in0(op_8_117__in0),
    .in1(op_8_117__in1),
    .out(op_8_117__out)
  );

  //Wire declarations for instance 'op_8_118' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_118__in0;
  wire [15:0] op_8_118__in1;
  wire [15:0] op_8_118__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_118(
    .in0(op_8_118__in0),
    .in1(op_8_118__in1),
    .out(op_8_118__out)
  );

  //Wire declarations for instance 'op_8_119' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_119__in0;
  wire [15:0] op_8_119__in1;
  wire [15:0] op_8_119__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_119(
    .in0(op_8_119__in0),
    .in1(op_8_119__in1),
    .out(op_8_119__out)
  );

  //Wire declarations for instance 'op_8_12' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_12__in0;
  wire [15:0] op_8_12__in1;
  wire [15:0] op_8_12__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_12(
    .in0(op_8_12__in0),
    .in1(op_8_12__in1),
    .out(op_8_12__out)
  );

  //Wire declarations for instance 'op_8_120' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_120__in0;
  wire [15:0] op_8_120__in1;
  wire [15:0] op_8_120__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_120(
    .in0(op_8_120__in0),
    .in1(op_8_120__in1),
    .out(op_8_120__out)
  );

  //Wire declarations for instance 'op_8_121' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_121__in0;
  wire [15:0] op_8_121__in1;
  wire [15:0] op_8_121__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_121(
    .in0(op_8_121__in0),
    .in1(op_8_121__in1),
    .out(op_8_121__out)
  );

  //Wire declarations for instance 'op_8_122' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_122__in0;
  wire [15:0] op_8_122__in1;
  wire [15:0] op_8_122__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_122(
    .in0(op_8_122__in0),
    .in1(op_8_122__in1),
    .out(op_8_122__out)
  );

  //Wire declarations for instance 'op_8_123' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_123__in0;
  wire [15:0] op_8_123__in1;
  wire [15:0] op_8_123__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_123(
    .in0(op_8_123__in0),
    .in1(op_8_123__in1),
    .out(op_8_123__out)
  );

  //Wire declarations for instance 'op_8_124' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_124__in0;
  wire [15:0] op_8_124__in1;
  wire [15:0] op_8_124__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_124(
    .in0(op_8_124__in0),
    .in1(op_8_124__in1),
    .out(op_8_124__out)
  );

  //Wire declarations for instance 'op_8_125' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_125__in0;
  wire [15:0] op_8_125__in1;
  wire [15:0] op_8_125__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_125(
    .in0(op_8_125__in0),
    .in1(op_8_125__in1),
    .out(op_8_125__out)
  );

  //Wire declarations for instance 'op_8_126' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_126__in0;
  wire [15:0] op_8_126__in1;
  wire [15:0] op_8_126__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_126(
    .in0(op_8_126__in0),
    .in1(op_8_126__in1),
    .out(op_8_126__out)
  );

  //Wire declarations for instance 'op_8_127' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_127__in0;
  wire [15:0] op_8_127__in1;
  wire [15:0] op_8_127__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_127(
    .in0(op_8_127__in0),
    .in1(op_8_127__in1),
    .out(op_8_127__out)
  );

  //Wire declarations for instance 'op_8_128' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_128__in0;
  wire [15:0] op_8_128__in1;
  wire [15:0] op_8_128__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_128(
    .in0(op_8_128__in0),
    .in1(op_8_128__in1),
    .out(op_8_128__out)
  );

  //Wire declarations for instance 'op_8_129' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_129__in0;
  wire [15:0] op_8_129__in1;
  wire [15:0] op_8_129__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_129(
    .in0(op_8_129__in0),
    .in1(op_8_129__in1),
    .out(op_8_129__out)
  );

  //Wire declarations for instance 'op_8_13' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_13__in0;
  wire [15:0] op_8_13__in1;
  wire [15:0] op_8_13__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_13(
    .in0(op_8_13__in0),
    .in1(op_8_13__in1),
    .out(op_8_13__out)
  );

  //Wire declarations for instance 'op_8_130' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_130__in0;
  wire [15:0] op_8_130__in1;
  wire [15:0] op_8_130__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_130(
    .in0(op_8_130__in0),
    .in1(op_8_130__in1),
    .out(op_8_130__out)
  );

  //Wire declarations for instance 'op_8_131' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_131__in0;
  wire [15:0] op_8_131__in1;
  wire [15:0] op_8_131__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_131(
    .in0(op_8_131__in0),
    .in1(op_8_131__in1),
    .out(op_8_131__out)
  );

  //Wire declarations for instance 'op_8_132' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_132__in0;
  wire [15:0] op_8_132__in1;
  wire [15:0] op_8_132__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_132(
    .in0(op_8_132__in0),
    .in1(op_8_132__in1),
    .out(op_8_132__out)
  );

  //Wire declarations for instance 'op_8_133' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_133__in0;
  wire [15:0] op_8_133__in1;
  wire [15:0] op_8_133__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_133(
    .in0(op_8_133__in0),
    .in1(op_8_133__in1),
    .out(op_8_133__out)
  );

  //Wire declarations for instance 'op_8_134' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_134__in0;
  wire [15:0] op_8_134__in1;
  wire [15:0] op_8_134__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_134(
    .in0(op_8_134__in0),
    .in1(op_8_134__in1),
    .out(op_8_134__out)
  );

  //Wire declarations for instance 'op_8_135' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_135__in0;
  wire [15:0] op_8_135__in1;
  wire [15:0] op_8_135__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_135(
    .in0(op_8_135__in0),
    .in1(op_8_135__in1),
    .out(op_8_135__out)
  );

  //Wire declarations for instance 'op_8_136' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_136__in0;
  wire [15:0] op_8_136__in1;
  wire [15:0] op_8_136__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_136(
    .in0(op_8_136__in0),
    .in1(op_8_136__in1),
    .out(op_8_136__out)
  );

  //Wire declarations for instance 'op_8_137' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_137__in0;
  wire [15:0] op_8_137__in1;
  wire [15:0] op_8_137__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_137(
    .in0(op_8_137__in0),
    .in1(op_8_137__in1),
    .out(op_8_137__out)
  );

  //Wire declarations for instance 'op_8_138' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_138__in0;
  wire [15:0] op_8_138__in1;
  wire [15:0] op_8_138__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_138(
    .in0(op_8_138__in0),
    .in1(op_8_138__in1),
    .out(op_8_138__out)
  );

  //Wire declarations for instance 'op_8_139' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_139__in0;
  wire [15:0] op_8_139__in1;
  wire [15:0] op_8_139__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_139(
    .in0(op_8_139__in0),
    .in1(op_8_139__in1),
    .out(op_8_139__out)
  );

  //Wire declarations for instance 'op_8_14' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_14__in0;
  wire [15:0] op_8_14__in1;
  wire [15:0] op_8_14__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_14(
    .in0(op_8_14__in0),
    .in1(op_8_14__in1),
    .out(op_8_14__out)
  );

  //Wire declarations for instance 'op_8_140' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_140__in0;
  wire [15:0] op_8_140__in1;
  wire [15:0] op_8_140__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_140(
    .in0(op_8_140__in0),
    .in1(op_8_140__in1),
    .out(op_8_140__out)
  );

  //Wire declarations for instance 'op_8_141' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_141__in0;
  wire [15:0] op_8_141__in1;
  wire [15:0] op_8_141__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_141(
    .in0(op_8_141__in0),
    .in1(op_8_141__in1),
    .out(op_8_141__out)
  );

  //Wire declarations for instance 'op_8_142' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_142__in0;
  wire [15:0] op_8_142__in1;
  wire [15:0] op_8_142__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_142(
    .in0(op_8_142__in0),
    .in1(op_8_142__in1),
    .out(op_8_142__out)
  );

  //Wire declarations for instance 'op_8_143' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_143__in0;
  wire [15:0] op_8_143__in1;
  wire [15:0] op_8_143__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_143(
    .in0(op_8_143__in0),
    .in1(op_8_143__in1),
    .out(op_8_143__out)
  );

  //Wire declarations for instance 'op_8_144' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_144__in0;
  wire [15:0] op_8_144__in1;
  wire [15:0] op_8_144__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_144(
    .in0(op_8_144__in0),
    .in1(op_8_144__in1),
    .out(op_8_144__out)
  );

  //Wire declarations for instance 'op_8_145' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_145__in0;
  wire [15:0] op_8_145__in1;
  wire [15:0] op_8_145__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_145(
    .in0(op_8_145__in0),
    .in1(op_8_145__in1),
    .out(op_8_145__out)
  );

  //Wire declarations for instance 'op_8_146' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_146__in0;
  wire [15:0] op_8_146__in1;
  wire [15:0] op_8_146__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_146(
    .in0(op_8_146__in0),
    .in1(op_8_146__in1),
    .out(op_8_146__out)
  );

  //Wire declarations for instance 'op_8_147' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_147__in0;
  wire [15:0] op_8_147__in1;
  wire [15:0] op_8_147__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_147(
    .in0(op_8_147__in0),
    .in1(op_8_147__in1),
    .out(op_8_147__out)
  );

  //Wire declarations for instance 'op_8_148' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_148__in0;
  wire [15:0] op_8_148__in1;
  wire [15:0] op_8_148__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_148(
    .in0(op_8_148__in0),
    .in1(op_8_148__in1),
    .out(op_8_148__out)
  );

  //Wire declarations for instance 'op_8_149' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_149__in0;
  wire [15:0] op_8_149__in1;
  wire [15:0] op_8_149__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_149(
    .in0(op_8_149__in0),
    .in1(op_8_149__in1),
    .out(op_8_149__out)
  );

  //Wire declarations for instance 'op_8_15' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_15__in0;
  wire [15:0] op_8_15__in1;
  wire [15:0] op_8_15__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_15(
    .in0(op_8_15__in0),
    .in1(op_8_15__in1),
    .out(op_8_15__out)
  );

  //Wire declarations for instance 'op_8_150' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_150__in0;
  wire [15:0] op_8_150__in1;
  wire [15:0] op_8_150__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_150(
    .in0(op_8_150__in0),
    .in1(op_8_150__in1),
    .out(op_8_150__out)
  );

  //Wire declarations for instance 'op_8_151' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_151__in0;
  wire [15:0] op_8_151__in1;
  wire [15:0] op_8_151__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_151(
    .in0(op_8_151__in0),
    .in1(op_8_151__in1),
    .out(op_8_151__out)
  );

  //Wire declarations for instance 'op_8_152' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_152__in0;
  wire [15:0] op_8_152__in1;
  wire [15:0] op_8_152__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_152(
    .in0(op_8_152__in0),
    .in1(op_8_152__in1),
    .out(op_8_152__out)
  );

  //Wire declarations for instance 'op_8_153' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_153__in0;
  wire [15:0] op_8_153__in1;
  wire [15:0] op_8_153__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_153(
    .in0(op_8_153__in0),
    .in1(op_8_153__in1),
    .out(op_8_153__out)
  );

  //Wire declarations for instance 'op_8_154' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_154__in0;
  wire [15:0] op_8_154__in1;
  wire [15:0] op_8_154__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_154(
    .in0(op_8_154__in0),
    .in1(op_8_154__in1),
    .out(op_8_154__out)
  );

  //Wire declarations for instance 'op_8_155' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_155__in0;
  wire [15:0] op_8_155__in1;
  wire [15:0] op_8_155__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_155(
    .in0(op_8_155__in0),
    .in1(op_8_155__in1),
    .out(op_8_155__out)
  );

  //Wire declarations for instance 'op_8_156' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_156__in0;
  wire [15:0] op_8_156__in1;
  wire [15:0] op_8_156__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_156(
    .in0(op_8_156__in0),
    .in1(op_8_156__in1),
    .out(op_8_156__out)
  );

  //Wire declarations for instance 'op_8_157' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_157__in0;
  wire [15:0] op_8_157__in1;
  wire [15:0] op_8_157__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_157(
    .in0(op_8_157__in0),
    .in1(op_8_157__in1),
    .out(op_8_157__out)
  );

  //Wire declarations for instance 'op_8_158' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_158__in0;
  wire [15:0] op_8_158__in1;
  wire [15:0] op_8_158__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_158(
    .in0(op_8_158__in0),
    .in1(op_8_158__in1),
    .out(op_8_158__out)
  );

  //Wire declarations for instance 'op_8_159' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_159__in0;
  wire [15:0] op_8_159__in1;
  wire [15:0] op_8_159__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_159(
    .in0(op_8_159__in0),
    .in1(op_8_159__in1),
    .out(op_8_159__out)
  );

  //Wire declarations for instance 'op_8_16' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_16__in0;
  wire [15:0] op_8_16__in1;
  wire [15:0] op_8_16__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_16(
    .in0(op_8_16__in0),
    .in1(op_8_16__in1),
    .out(op_8_16__out)
  );

  //Wire declarations for instance 'op_8_160' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_160__in0;
  wire [15:0] op_8_160__in1;
  wire [15:0] op_8_160__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_160(
    .in0(op_8_160__in0),
    .in1(op_8_160__in1),
    .out(op_8_160__out)
  );

  //Wire declarations for instance 'op_8_161' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_161__in0;
  wire [15:0] op_8_161__in1;
  wire [15:0] op_8_161__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_161(
    .in0(op_8_161__in0),
    .in1(op_8_161__in1),
    .out(op_8_161__out)
  );

  //Wire declarations for instance 'op_8_162' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_162__in0;
  wire [15:0] op_8_162__in1;
  wire [15:0] op_8_162__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_162(
    .in0(op_8_162__in0),
    .in1(op_8_162__in1),
    .out(op_8_162__out)
  );

  //Wire declarations for instance 'op_8_163' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_163__in0;
  wire [15:0] op_8_163__in1;
  wire [15:0] op_8_163__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_163(
    .in0(op_8_163__in0),
    .in1(op_8_163__in1),
    .out(op_8_163__out)
  );

  //Wire declarations for instance 'op_8_164' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_164__in0;
  wire [15:0] op_8_164__in1;
  wire [15:0] op_8_164__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_164(
    .in0(op_8_164__in0),
    .in1(op_8_164__in1),
    .out(op_8_164__out)
  );

  //Wire declarations for instance 'op_8_165' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_165__in0;
  wire [15:0] op_8_165__in1;
  wire [15:0] op_8_165__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_165(
    .in0(op_8_165__in0),
    .in1(op_8_165__in1),
    .out(op_8_165__out)
  );

  //Wire declarations for instance 'op_8_166' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_166__in0;
  wire [15:0] op_8_166__in1;
  wire [15:0] op_8_166__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_166(
    .in0(op_8_166__in0),
    .in1(op_8_166__in1),
    .out(op_8_166__out)
  );

  //Wire declarations for instance 'op_8_167' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_167__in0;
  wire [15:0] op_8_167__in1;
  wire [15:0] op_8_167__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_167(
    .in0(op_8_167__in0),
    .in1(op_8_167__in1),
    .out(op_8_167__out)
  );

  //Wire declarations for instance 'op_8_168' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_168__in0;
  wire [15:0] op_8_168__in1;
  wire [15:0] op_8_168__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_168(
    .in0(op_8_168__in0),
    .in1(op_8_168__in1),
    .out(op_8_168__out)
  );

  //Wire declarations for instance 'op_8_169' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_169__in0;
  wire [15:0] op_8_169__in1;
  wire [15:0] op_8_169__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_169(
    .in0(op_8_169__in0),
    .in1(op_8_169__in1),
    .out(op_8_169__out)
  );

  //Wire declarations for instance 'op_8_17' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_17__in0;
  wire [15:0] op_8_17__in1;
  wire [15:0] op_8_17__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_17(
    .in0(op_8_17__in0),
    .in1(op_8_17__in1),
    .out(op_8_17__out)
  );

  //Wire declarations for instance 'op_8_170' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_170__in0;
  wire [15:0] op_8_170__in1;
  wire [15:0] op_8_170__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_170(
    .in0(op_8_170__in0),
    .in1(op_8_170__in1),
    .out(op_8_170__out)
  );

  //Wire declarations for instance 'op_8_171' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_171__in0;
  wire [15:0] op_8_171__in1;
  wire [15:0] op_8_171__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_171(
    .in0(op_8_171__in0),
    .in1(op_8_171__in1),
    .out(op_8_171__out)
  );

  //Wire declarations for instance 'op_8_172' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_172__in0;
  wire [15:0] op_8_172__in1;
  wire [15:0] op_8_172__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_172(
    .in0(op_8_172__in0),
    .in1(op_8_172__in1),
    .out(op_8_172__out)
  );

  //Wire declarations for instance 'op_8_173' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_173__in0;
  wire [15:0] op_8_173__in1;
  wire [15:0] op_8_173__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_173(
    .in0(op_8_173__in0),
    .in1(op_8_173__in1),
    .out(op_8_173__out)
  );

  //Wire declarations for instance 'op_8_174' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_174__in0;
  wire [15:0] op_8_174__in1;
  wire [15:0] op_8_174__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_174(
    .in0(op_8_174__in0),
    .in1(op_8_174__in1),
    .out(op_8_174__out)
  );

  //Wire declarations for instance 'op_8_175' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_175__in0;
  wire [15:0] op_8_175__in1;
  wire [15:0] op_8_175__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_175(
    .in0(op_8_175__in0),
    .in1(op_8_175__in1),
    .out(op_8_175__out)
  );

  //Wire declarations for instance 'op_8_176' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_176__in0;
  wire [15:0] op_8_176__in1;
  wire [15:0] op_8_176__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_176(
    .in0(op_8_176__in0),
    .in1(op_8_176__in1),
    .out(op_8_176__out)
  );

  //Wire declarations for instance 'op_8_177' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_177__in0;
  wire [15:0] op_8_177__in1;
  wire [15:0] op_8_177__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_177(
    .in0(op_8_177__in0),
    .in1(op_8_177__in1),
    .out(op_8_177__out)
  );

  //Wire declarations for instance 'op_8_178' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_178__in0;
  wire [15:0] op_8_178__in1;
  wire [15:0] op_8_178__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_178(
    .in0(op_8_178__in0),
    .in1(op_8_178__in1),
    .out(op_8_178__out)
  );

  //Wire declarations for instance 'op_8_179' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_179__in0;
  wire [15:0] op_8_179__in1;
  wire [15:0] op_8_179__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_179(
    .in0(op_8_179__in0),
    .in1(op_8_179__in1),
    .out(op_8_179__out)
  );

  //Wire declarations for instance 'op_8_18' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_18__in0;
  wire [15:0] op_8_18__in1;
  wire [15:0] op_8_18__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_18(
    .in0(op_8_18__in0),
    .in1(op_8_18__in1),
    .out(op_8_18__out)
  );

  //Wire declarations for instance 'op_8_180' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_180__in0;
  wire [15:0] op_8_180__in1;
  wire [15:0] op_8_180__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_180(
    .in0(op_8_180__in0),
    .in1(op_8_180__in1),
    .out(op_8_180__out)
  );

  //Wire declarations for instance 'op_8_181' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_181__in0;
  wire [15:0] op_8_181__in1;
  wire [15:0] op_8_181__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_181(
    .in0(op_8_181__in0),
    .in1(op_8_181__in1),
    .out(op_8_181__out)
  );

  //Wire declarations for instance 'op_8_182' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_182__in0;
  wire [15:0] op_8_182__in1;
  wire [15:0] op_8_182__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_182(
    .in0(op_8_182__in0),
    .in1(op_8_182__in1),
    .out(op_8_182__out)
  );

  //Wire declarations for instance 'op_8_183' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_183__in0;
  wire [15:0] op_8_183__in1;
  wire [15:0] op_8_183__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_183(
    .in0(op_8_183__in0),
    .in1(op_8_183__in1),
    .out(op_8_183__out)
  );

  //Wire declarations for instance 'op_8_184' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_184__in0;
  wire [15:0] op_8_184__in1;
  wire [15:0] op_8_184__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_184(
    .in0(op_8_184__in0),
    .in1(op_8_184__in1),
    .out(op_8_184__out)
  );

  //Wire declarations for instance 'op_8_185' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_185__in0;
  wire [15:0] op_8_185__in1;
  wire [15:0] op_8_185__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_185(
    .in0(op_8_185__in0),
    .in1(op_8_185__in1),
    .out(op_8_185__out)
  );

  //Wire declarations for instance 'op_8_186' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_186__in0;
  wire [15:0] op_8_186__in1;
  wire [15:0] op_8_186__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_186(
    .in0(op_8_186__in0),
    .in1(op_8_186__in1),
    .out(op_8_186__out)
  );

  //Wire declarations for instance 'op_8_187' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_187__in0;
  wire [15:0] op_8_187__in1;
  wire [15:0] op_8_187__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_187(
    .in0(op_8_187__in0),
    .in1(op_8_187__in1),
    .out(op_8_187__out)
  );

  //Wire declarations for instance 'op_8_188' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_188__in0;
  wire [15:0] op_8_188__in1;
  wire [15:0] op_8_188__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_188(
    .in0(op_8_188__in0),
    .in1(op_8_188__in1),
    .out(op_8_188__out)
  );

  //Wire declarations for instance 'op_8_189' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_189__in0;
  wire [15:0] op_8_189__in1;
  wire [15:0] op_8_189__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_189(
    .in0(op_8_189__in0),
    .in1(op_8_189__in1),
    .out(op_8_189__out)
  );

  //Wire declarations for instance 'op_8_19' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_19__in0;
  wire [15:0] op_8_19__in1;
  wire [15:0] op_8_19__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_19(
    .in0(op_8_19__in0),
    .in1(op_8_19__in1),
    .out(op_8_19__out)
  );

  //Wire declarations for instance 'op_8_190' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_190__in0;
  wire [15:0] op_8_190__in1;
  wire [15:0] op_8_190__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_190(
    .in0(op_8_190__in0),
    .in1(op_8_190__in1),
    .out(op_8_190__out)
  );

  //Wire declarations for instance 'op_8_191' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_191__in0;
  wire [15:0] op_8_191__in1;
  wire [15:0] op_8_191__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_191(
    .in0(op_8_191__in0),
    .in1(op_8_191__in1),
    .out(op_8_191__out)
  );

  //Wire declarations for instance 'op_8_192' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_192__in0;
  wire [15:0] op_8_192__in1;
  wire [15:0] op_8_192__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_192(
    .in0(op_8_192__in0),
    .in1(op_8_192__in1),
    .out(op_8_192__out)
  );

  //Wire declarations for instance 'op_8_193' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_193__in0;
  wire [15:0] op_8_193__in1;
  wire [15:0] op_8_193__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_193(
    .in0(op_8_193__in0),
    .in1(op_8_193__in1),
    .out(op_8_193__out)
  );

  //Wire declarations for instance 'op_8_194' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_194__in0;
  wire [15:0] op_8_194__in1;
  wire [15:0] op_8_194__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_194(
    .in0(op_8_194__in0),
    .in1(op_8_194__in1),
    .out(op_8_194__out)
  );

  //Wire declarations for instance 'op_8_195' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_195__in0;
  wire [15:0] op_8_195__in1;
  wire [15:0] op_8_195__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_195(
    .in0(op_8_195__in0),
    .in1(op_8_195__in1),
    .out(op_8_195__out)
  );

  //Wire declarations for instance 'op_8_196' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_196__in0;
  wire [15:0] op_8_196__in1;
  wire [15:0] op_8_196__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_196(
    .in0(op_8_196__in0),
    .in1(op_8_196__in1),
    .out(op_8_196__out)
  );

  //Wire declarations for instance 'op_8_197' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_197__in0;
  wire [15:0] op_8_197__in1;
  wire [15:0] op_8_197__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_197(
    .in0(op_8_197__in0),
    .in1(op_8_197__in1),
    .out(op_8_197__out)
  );

  //Wire declarations for instance 'op_8_198' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_198__in0;
  wire [15:0] op_8_198__in1;
  wire [15:0] op_8_198__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_198(
    .in0(op_8_198__in0),
    .in1(op_8_198__in1),
    .out(op_8_198__out)
  );

  //Wire declarations for instance 'op_8_199' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_199__in0;
  wire [15:0] op_8_199__in1;
  wire [15:0] op_8_199__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_199(
    .in0(op_8_199__in0),
    .in1(op_8_199__in1),
    .out(op_8_199__out)
  );

  //Wire declarations for instance 'op_8_2' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_2__in0;
  wire [15:0] op_8_2__in1;
  wire [15:0] op_8_2__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_2(
    .in0(op_8_2__in0),
    .in1(op_8_2__in1),
    .out(op_8_2__out)
  );

  //Wire declarations for instance 'op_8_20' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_20__in0;
  wire [15:0] op_8_20__in1;
  wire [15:0] op_8_20__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_20(
    .in0(op_8_20__in0),
    .in1(op_8_20__in1),
    .out(op_8_20__out)
  );

  //Wire declarations for instance 'op_8_200' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_200__in0;
  wire [15:0] op_8_200__in1;
  wire [15:0] op_8_200__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_200(
    .in0(op_8_200__in0),
    .in1(op_8_200__in1),
    .out(op_8_200__out)
  );

  //Wire declarations for instance 'op_8_201' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_201__in0;
  wire [15:0] op_8_201__in1;
  wire [15:0] op_8_201__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_201(
    .in0(op_8_201__in0),
    .in1(op_8_201__in1),
    .out(op_8_201__out)
  );

  //Wire declarations for instance 'op_8_202' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_202__in0;
  wire [15:0] op_8_202__in1;
  wire [15:0] op_8_202__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_202(
    .in0(op_8_202__in0),
    .in1(op_8_202__in1),
    .out(op_8_202__out)
  );

  //Wire declarations for instance 'op_8_203' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_203__in0;
  wire [15:0] op_8_203__in1;
  wire [15:0] op_8_203__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_203(
    .in0(op_8_203__in0),
    .in1(op_8_203__in1),
    .out(op_8_203__out)
  );

  //Wire declarations for instance 'op_8_204' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_204__in0;
  wire [15:0] op_8_204__in1;
  wire [15:0] op_8_204__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_204(
    .in0(op_8_204__in0),
    .in1(op_8_204__in1),
    .out(op_8_204__out)
  );

  //Wire declarations for instance 'op_8_205' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_205__in0;
  wire [15:0] op_8_205__in1;
  wire [15:0] op_8_205__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_205(
    .in0(op_8_205__in0),
    .in1(op_8_205__in1),
    .out(op_8_205__out)
  );

  //Wire declarations for instance 'op_8_206' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_206__in0;
  wire [15:0] op_8_206__in1;
  wire [15:0] op_8_206__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_206(
    .in0(op_8_206__in0),
    .in1(op_8_206__in1),
    .out(op_8_206__out)
  );

  //Wire declarations for instance 'op_8_207' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_207__in0;
  wire [15:0] op_8_207__in1;
  wire [15:0] op_8_207__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_207(
    .in0(op_8_207__in0),
    .in1(op_8_207__in1),
    .out(op_8_207__out)
  );

  //Wire declarations for instance 'op_8_208' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_208__in0;
  wire [15:0] op_8_208__in1;
  wire [15:0] op_8_208__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_208(
    .in0(op_8_208__in0),
    .in1(op_8_208__in1),
    .out(op_8_208__out)
  );

  //Wire declarations for instance 'op_8_209' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_209__in0;
  wire [15:0] op_8_209__in1;
  wire [15:0] op_8_209__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_209(
    .in0(op_8_209__in0),
    .in1(op_8_209__in1),
    .out(op_8_209__out)
  );

  //Wire declarations for instance 'op_8_21' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_21__in0;
  wire [15:0] op_8_21__in1;
  wire [15:0] op_8_21__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_21(
    .in0(op_8_21__in0),
    .in1(op_8_21__in1),
    .out(op_8_21__out)
  );

  //Wire declarations for instance 'op_8_210' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_210__in0;
  wire [15:0] op_8_210__in1;
  wire [15:0] op_8_210__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_210(
    .in0(op_8_210__in0),
    .in1(op_8_210__in1),
    .out(op_8_210__out)
  );

  //Wire declarations for instance 'op_8_211' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_211__in0;
  wire [15:0] op_8_211__in1;
  wire [15:0] op_8_211__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_211(
    .in0(op_8_211__in0),
    .in1(op_8_211__in1),
    .out(op_8_211__out)
  );

  //Wire declarations for instance 'op_8_212' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_212__in0;
  wire [15:0] op_8_212__in1;
  wire [15:0] op_8_212__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_212(
    .in0(op_8_212__in0),
    .in1(op_8_212__in1),
    .out(op_8_212__out)
  );

  //Wire declarations for instance 'op_8_213' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_213__in0;
  wire [15:0] op_8_213__in1;
  wire [15:0] op_8_213__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_213(
    .in0(op_8_213__in0),
    .in1(op_8_213__in1),
    .out(op_8_213__out)
  );

  //Wire declarations for instance 'op_8_214' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_214__in0;
  wire [15:0] op_8_214__in1;
  wire [15:0] op_8_214__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_214(
    .in0(op_8_214__in0),
    .in1(op_8_214__in1),
    .out(op_8_214__out)
  );

  //Wire declarations for instance 'op_8_215' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_215__in0;
  wire [15:0] op_8_215__in1;
  wire [15:0] op_8_215__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_215(
    .in0(op_8_215__in0),
    .in1(op_8_215__in1),
    .out(op_8_215__out)
  );

  //Wire declarations for instance 'op_8_216' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_216__in0;
  wire [15:0] op_8_216__in1;
  wire [15:0] op_8_216__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_216(
    .in0(op_8_216__in0),
    .in1(op_8_216__in1),
    .out(op_8_216__out)
  );

  //Wire declarations for instance 'op_8_217' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_217__in0;
  wire [15:0] op_8_217__in1;
  wire [15:0] op_8_217__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_217(
    .in0(op_8_217__in0),
    .in1(op_8_217__in1),
    .out(op_8_217__out)
  );

  //Wire declarations for instance 'op_8_218' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_218__in0;
  wire [15:0] op_8_218__in1;
  wire [15:0] op_8_218__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_218(
    .in0(op_8_218__in0),
    .in1(op_8_218__in1),
    .out(op_8_218__out)
  );

  //Wire declarations for instance 'op_8_219' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_219__in0;
  wire [15:0] op_8_219__in1;
  wire [15:0] op_8_219__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_219(
    .in0(op_8_219__in0),
    .in1(op_8_219__in1),
    .out(op_8_219__out)
  );

  //Wire declarations for instance 'op_8_22' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_22__in0;
  wire [15:0] op_8_22__in1;
  wire [15:0] op_8_22__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_22(
    .in0(op_8_22__in0),
    .in1(op_8_22__in1),
    .out(op_8_22__out)
  );

  //Wire declarations for instance 'op_8_220' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_220__in0;
  wire [15:0] op_8_220__in1;
  wire [15:0] op_8_220__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_220(
    .in0(op_8_220__in0),
    .in1(op_8_220__in1),
    .out(op_8_220__out)
  );

  //Wire declarations for instance 'op_8_221' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_221__in0;
  wire [15:0] op_8_221__in1;
  wire [15:0] op_8_221__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_221(
    .in0(op_8_221__in0),
    .in1(op_8_221__in1),
    .out(op_8_221__out)
  );

  //Wire declarations for instance 'op_8_222' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_222__in0;
  wire [15:0] op_8_222__in1;
  wire [15:0] op_8_222__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_222(
    .in0(op_8_222__in0),
    .in1(op_8_222__in1),
    .out(op_8_222__out)
  );

  //Wire declarations for instance 'op_8_223' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_223__in0;
  wire [15:0] op_8_223__in1;
  wire [15:0] op_8_223__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_223(
    .in0(op_8_223__in0),
    .in1(op_8_223__in1),
    .out(op_8_223__out)
  );

  //Wire declarations for instance 'op_8_224' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_224__in0;
  wire [15:0] op_8_224__in1;
  wire [15:0] op_8_224__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_224(
    .in0(op_8_224__in0),
    .in1(op_8_224__in1),
    .out(op_8_224__out)
  );

  //Wire declarations for instance 'op_8_225' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_225__in0;
  wire [15:0] op_8_225__in1;
  wire [15:0] op_8_225__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_225(
    .in0(op_8_225__in0),
    .in1(op_8_225__in1),
    .out(op_8_225__out)
  );

  //Wire declarations for instance 'op_8_226' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_226__in0;
  wire [15:0] op_8_226__in1;
  wire [15:0] op_8_226__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_226(
    .in0(op_8_226__in0),
    .in1(op_8_226__in1),
    .out(op_8_226__out)
  );

  //Wire declarations for instance 'op_8_227' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_227__in0;
  wire [15:0] op_8_227__in1;
  wire [15:0] op_8_227__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_227(
    .in0(op_8_227__in0),
    .in1(op_8_227__in1),
    .out(op_8_227__out)
  );

  //Wire declarations for instance 'op_8_228' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_228__in0;
  wire [15:0] op_8_228__in1;
  wire [15:0] op_8_228__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_228(
    .in0(op_8_228__in0),
    .in1(op_8_228__in1),
    .out(op_8_228__out)
  );

  //Wire declarations for instance 'op_8_229' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_229__in0;
  wire [15:0] op_8_229__in1;
  wire [15:0] op_8_229__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_229(
    .in0(op_8_229__in0),
    .in1(op_8_229__in1),
    .out(op_8_229__out)
  );

  //Wire declarations for instance 'op_8_23' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_23__in0;
  wire [15:0] op_8_23__in1;
  wire [15:0] op_8_23__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_23(
    .in0(op_8_23__in0),
    .in1(op_8_23__in1),
    .out(op_8_23__out)
  );

  //Wire declarations for instance 'op_8_230' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_230__in0;
  wire [15:0] op_8_230__in1;
  wire [15:0] op_8_230__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_230(
    .in0(op_8_230__in0),
    .in1(op_8_230__in1),
    .out(op_8_230__out)
  );

  //Wire declarations for instance 'op_8_231' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_231__in0;
  wire [15:0] op_8_231__in1;
  wire [15:0] op_8_231__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_231(
    .in0(op_8_231__in0),
    .in1(op_8_231__in1),
    .out(op_8_231__out)
  );

  //Wire declarations for instance 'op_8_232' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_232__in0;
  wire [15:0] op_8_232__in1;
  wire [15:0] op_8_232__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_232(
    .in0(op_8_232__in0),
    .in1(op_8_232__in1),
    .out(op_8_232__out)
  );

  //Wire declarations for instance 'op_8_233' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_233__in0;
  wire [15:0] op_8_233__in1;
  wire [15:0] op_8_233__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_233(
    .in0(op_8_233__in0),
    .in1(op_8_233__in1),
    .out(op_8_233__out)
  );

  //Wire declarations for instance 'op_8_234' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_234__in0;
  wire [15:0] op_8_234__in1;
  wire [15:0] op_8_234__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_234(
    .in0(op_8_234__in0),
    .in1(op_8_234__in1),
    .out(op_8_234__out)
  );

  //Wire declarations for instance 'op_8_235' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_235__in0;
  wire [15:0] op_8_235__in1;
  wire [15:0] op_8_235__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_235(
    .in0(op_8_235__in0),
    .in1(op_8_235__in1),
    .out(op_8_235__out)
  );

  //Wire declarations for instance 'op_8_236' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_236__in0;
  wire [15:0] op_8_236__in1;
  wire [15:0] op_8_236__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_236(
    .in0(op_8_236__in0),
    .in1(op_8_236__in1),
    .out(op_8_236__out)
  );

  //Wire declarations for instance 'op_8_237' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_237__in0;
  wire [15:0] op_8_237__in1;
  wire [15:0] op_8_237__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_237(
    .in0(op_8_237__in0),
    .in1(op_8_237__in1),
    .out(op_8_237__out)
  );

  //Wire declarations for instance 'op_8_238' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_238__in0;
  wire [15:0] op_8_238__in1;
  wire [15:0] op_8_238__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_238(
    .in0(op_8_238__in0),
    .in1(op_8_238__in1),
    .out(op_8_238__out)
  );

  //Wire declarations for instance 'op_8_239' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_239__in0;
  wire [15:0] op_8_239__in1;
  wire [15:0] op_8_239__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_239(
    .in0(op_8_239__in0),
    .in1(op_8_239__in1),
    .out(op_8_239__out)
  );

  //Wire declarations for instance 'op_8_24' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_24__in0;
  wire [15:0] op_8_24__in1;
  wire [15:0] op_8_24__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_24(
    .in0(op_8_24__in0),
    .in1(op_8_24__in1),
    .out(op_8_24__out)
  );

  //Wire declarations for instance 'op_8_240' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_240__in0;
  wire [15:0] op_8_240__in1;
  wire [15:0] op_8_240__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_240(
    .in0(op_8_240__in0),
    .in1(op_8_240__in1),
    .out(op_8_240__out)
  );

  //Wire declarations for instance 'op_8_241' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_241__in0;
  wire [15:0] op_8_241__in1;
  wire [15:0] op_8_241__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_241(
    .in0(op_8_241__in0),
    .in1(op_8_241__in1),
    .out(op_8_241__out)
  );

  //Wire declarations for instance 'op_8_242' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_242__in0;
  wire [15:0] op_8_242__in1;
  wire [15:0] op_8_242__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_242(
    .in0(op_8_242__in0),
    .in1(op_8_242__in1),
    .out(op_8_242__out)
  );

  //Wire declarations for instance 'op_8_243' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_243__in0;
  wire [15:0] op_8_243__in1;
  wire [15:0] op_8_243__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_243(
    .in0(op_8_243__in0),
    .in1(op_8_243__in1),
    .out(op_8_243__out)
  );

  //Wire declarations for instance 'op_8_244' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_244__in0;
  wire [15:0] op_8_244__in1;
  wire [15:0] op_8_244__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_244(
    .in0(op_8_244__in0),
    .in1(op_8_244__in1),
    .out(op_8_244__out)
  );

  //Wire declarations for instance 'op_8_245' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_245__in0;
  wire [15:0] op_8_245__in1;
  wire [15:0] op_8_245__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_245(
    .in0(op_8_245__in0),
    .in1(op_8_245__in1),
    .out(op_8_245__out)
  );

  //Wire declarations for instance 'op_8_246' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_246__in0;
  wire [15:0] op_8_246__in1;
  wire [15:0] op_8_246__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_246(
    .in0(op_8_246__in0),
    .in1(op_8_246__in1),
    .out(op_8_246__out)
  );

  //Wire declarations for instance 'op_8_247' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_247__in0;
  wire [15:0] op_8_247__in1;
  wire [15:0] op_8_247__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_247(
    .in0(op_8_247__in0),
    .in1(op_8_247__in1),
    .out(op_8_247__out)
  );

  //Wire declarations for instance 'op_8_248' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_248__in0;
  wire [15:0] op_8_248__in1;
  wire [15:0] op_8_248__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_248(
    .in0(op_8_248__in0),
    .in1(op_8_248__in1),
    .out(op_8_248__out)
  );

  //Wire declarations for instance 'op_8_249' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_249__in0;
  wire [15:0] op_8_249__in1;
  wire [15:0] op_8_249__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_249(
    .in0(op_8_249__in0),
    .in1(op_8_249__in1),
    .out(op_8_249__out)
  );

  //Wire declarations for instance 'op_8_25' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_25__in0;
  wire [15:0] op_8_25__in1;
  wire [15:0] op_8_25__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_25(
    .in0(op_8_25__in0),
    .in1(op_8_25__in1),
    .out(op_8_25__out)
  );

  //Wire declarations for instance 'op_8_250' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_250__in0;
  wire [15:0] op_8_250__in1;
  wire [15:0] op_8_250__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_250(
    .in0(op_8_250__in0),
    .in1(op_8_250__in1),
    .out(op_8_250__out)
  );

  //Wire declarations for instance 'op_8_251' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_251__in0;
  wire [15:0] op_8_251__in1;
  wire [15:0] op_8_251__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_251(
    .in0(op_8_251__in0),
    .in1(op_8_251__in1),
    .out(op_8_251__out)
  );

  //Wire declarations for instance 'op_8_252' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_252__in0;
  wire [15:0] op_8_252__in1;
  wire [15:0] op_8_252__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_252(
    .in0(op_8_252__in0),
    .in1(op_8_252__in1),
    .out(op_8_252__out)
  );

  //Wire declarations for instance 'op_8_253' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_253__in0;
  wire [15:0] op_8_253__in1;
  wire [15:0] op_8_253__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_253(
    .in0(op_8_253__in0),
    .in1(op_8_253__in1),
    .out(op_8_253__out)
  );

  //Wire declarations for instance 'op_8_254' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_254__in0;
  wire [15:0] op_8_254__in1;
  wire [15:0] op_8_254__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_254(
    .in0(op_8_254__in0),
    .in1(op_8_254__in1),
    .out(op_8_254__out)
  );

  //Wire declarations for instance 'op_8_255' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_255__in0;
  wire [15:0] op_8_255__in1;
  wire [15:0] op_8_255__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_255(
    .in0(op_8_255__in0),
    .in1(op_8_255__in1),
    .out(op_8_255__out)
  );

  //Wire declarations for instance 'op_8_26' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_26__in0;
  wire [15:0] op_8_26__in1;
  wire [15:0] op_8_26__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_26(
    .in0(op_8_26__in0),
    .in1(op_8_26__in1),
    .out(op_8_26__out)
  );

  //Wire declarations for instance 'op_8_27' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_27__in0;
  wire [15:0] op_8_27__in1;
  wire [15:0] op_8_27__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_27(
    .in0(op_8_27__in0),
    .in1(op_8_27__in1),
    .out(op_8_27__out)
  );

  //Wire declarations for instance 'op_8_28' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_28__in0;
  wire [15:0] op_8_28__in1;
  wire [15:0] op_8_28__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_28(
    .in0(op_8_28__in0),
    .in1(op_8_28__in1),
    .out(op_8_28__out)
  );

  //Wire declarations for instance 'op_8_29' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_29__in0;
  wire [15:0] op_8_29__in1;
  wire [15:0] op_8_29__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_29(
    .in0(op_8_29__in0),
    .in1(op_8_29__in1),
    .out(op_8_29__out)
  );

  //Wire declarations for instance 'op_8_3' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_3__in0;
  wire [15:0] op_8_3__in1;
  wire [15:0] op_8_3__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_3(
    .in0(op_8_3__in0),
    .in1(op_8_3__in1),
    .out(op_8_3__out)
  );

  //Wire declarations for instance 'op_8_30' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_30__in0;
  wire [15:0] op_8_30__in1;
  wire [15:0] op_8_30__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_30(
    .in0(op_8_30__in0),
    .in1(op_8_30__in1),
    .out(op_8_30__out)
  );

  //Wire declarations for instance 'op_8_31' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_31__in0;
  wire [15:0] op_8_31__in1;
  wire [15:0] op_8_31__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_31(
    .in0(op_8_31__in0),
    .in1(op_8_31__in1),
    .out(op_8_31__out)
  );

  //Wire declarations for instance 'op_8_32' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_32__in0;
  wire [15:0] op_8_32__in1;
  wire [15:0] op_8_32__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_32(
    .in0(op_8_32__in0),
    .in1(op_8_32__in1),
    .out(op_8_32__out)
  );

  //Wire declarations for instance 'op_8_33' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_33__in0;
  wire [15:0] op_8_33__in1;
  wire [15:0] op_8_33__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_33(
    .in0(op_8_33__in0),
    .in1(op_8_33__in1),
    .out(op_8_33__out)
  );

  //Wire declarations for instance 'op_8_34' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_34__in0;
  wire [15:0] op_8_34__in1;
  wire [15:0] op_8_34__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_34(
    .in0(op_8_34__in0),
    .in1(op_8_34__in1),
    .out(op_8_34__out)
  );

  //Wire declarations for instance 'op_8_35' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_35__in0;
  wire [15:0] op_8_35__in1;
  wire [15:0] op_8_35__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_35(
    .in0(op_8_35__in0),
    .in1(op_8_35__in1),
    .out(op_8_35__out)
  );

  //Wire declarations for instance 'op_8_36' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_36__in0;
  wire [15:0] op_8_36__in1;
  wire [15:0] op_8_36__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_36(
    .in0(op_8_36__in0),
    .in1(op_8_36__in1),
    .out(op_8_36__out)
  );

  //Wire declarations for instance 'op_8_37' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_37__in0;
  wire [15:0] op_8_37__in1;
  wire [15:0] op_8_37__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_37(
    .in0(op_8_37__in0),
    .in1(op_8_37__in1),
    .out(op_8_37__out)
  );

  //Wire declarations for instance 'op_8_38' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_38__in0;
  wire [15:0] op_8_38__in1;
  wire [15:0] op_8_38__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_38(
    .in0(op_8_38__in0),
    .in1(op_8_38__in1),
    .out(op_8_38__out)
  );

  //Wire declarations for instance 'op_8_39' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_39__in0;
  wire [15:0] op_8_39__in1;
  wire [15:0] op_8_39__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_39(
    .in0(op_8_39__in0),
    .in1(op_8_39__in1),
    .out(op_8_39__out)
  );

  //Wire declarations for instance 'op_8_4' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_4__in0;
  wire [15:0] op_8_4__in1;
  wire [15:0] op_8_4__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_4(
    .in0(op_8_4__in0),
    .in1(op_8_4__in1),
    .out(op_8_4__out)
  );

  //Wire declarations for instance 'op_8_40' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_40__in0;
  wire [15:0] op_8_40__in1;
  wire [15:0] op_8_40__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_40(
    .in0(op_8_40__in0),
    .in1(op_8_40__in1),
    .out(op_8_40__out)
  );

  //Wire declarations for instance 'op_8_41' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_41__in0;
  wire [15:0] op_8_41__in1;
  wire [15:0] op_8_41__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_41(
    .in0(op_8_41__in0),
    .in1(op_8_41__in1),
    .out(op_8_41__out)
  );

  //Wire declarations for instance 'op_8_42' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_42__in0;
  wire [15:0] op_8_42__in1;
  wire [15:0] op_8_42__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_42(
    .in0(op_8_42__in0),
    .in1(op_8_42__in1),
    .out(op_8_42__out)
  );

  //Wire declarations for instance 'op_8_43' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_43__in0;
  wire [15:0] op_8_43__in1;
  wire [15:0] op_8_43__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_43(
    .in0(op_8_43__in0),
    .in1(op_8_43__in1),
    .out(op_8_43__out)
  );

  //Wire declarations for instance 'op_8_44' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_44__in0;
  wire [15:0] op_8_44__in1;
  wire [15:0] op_8_44__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_44(
    .in0(op_8_44__in0),
    .in1(op_8_44__in1),
    .out(op_8_44__out)
  );

  //Wire declarations for instance 'op_8_45' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_45__in0;
  wire [15:0] op_8_45__in1;
  wire [15:0] op_8_45__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_45(
    .in0(op_8_45__in0),
    .in1(op_8_45__in1),
    .out(op_8_45__out)
  );

  //Wire declarations for instance 'op_8_46' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_46__in0;
  wire [15:0] op_8_46__in1;
  wire [15:0] op_8_46__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_46(
    .in0(op_8_46__in0),
    .in1(op_8_46__in1),
    .out(op_8_46__out)
  );

  //Wire declarations for instance 'op_8_47' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_47__in0;
  wire [15:0] op_8_47__in1;
  wire [15:0] op_8_47__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_47(
    .in0(op_8_47__in0),
    .in1(op_8_47__in1),
    .out(op_8_47__out)
  );

  //Wire declarations for instance 'op_8_48' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_48__in0;
  wire [15:0] op_8_48__in1;
  wire [15:0] op_8_48__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_48(
    .in0(op_8_48__in0),
    .in1(op_8_48__in1),
    .out(op_8_48__out)
  );

  //Wire declarations for instance 'op_8_49' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_49__in0;
  wire [15:0] op_8_49__in1;
  wire [15:0] op_8_49__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_49(
    .in0(op_8_49__in0),
    .in1(op_8_49__in1),
    .out(op_8_49__out)
  );

  //Wire declarations for instance 'op_8_5' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_5__in0;
  wire [15:0] op_8_5__in1;
  wire [15:0] op_8_5__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_5(
    .in0(op_8_5__in0),
    .in1(op_8_5__in1),
    .out(op_8_5__out)
  );

  //Wire declarations for instance 'op_8_50' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_50__in0;
  wire [15:0] op_8_50__in1;
  wire [15:0] op_8_50__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_50(
    .in0(op_8_50__in0),
    .in1(op_8_50__in1),
    .out(op_8_50__out)
  );

  //Wire declarations for instance 'op_8_51' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_51__in0;
  wire [15:0] op_8_51__in1;
  wire [15:0] op_8_51__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_51(
    .in0(op_8_51__in0),
    .in1(op_8_51__in1),
    .out(op_8_51__out)
  );

  //Wire declarations for instance 'op_8_52' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_52__in0;
  wire [15:0] op_8_52__in1;
  wire [15:0] op_8_52__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_52(
    .in0(op_8_52__in0),
    .in1(op_8_52__in1),
    .out(op_8_52__out)
  );

  //Wire declarations for instance 'op_8_53' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_53__in0;
  wire [15:0] op_8_53__in1;
  wire [15:0] op_8_53__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_53(
    .in0(op_8_53__in0),
    .in1(op_8_53__in1),
    .out(op_8_53__out)
  );

  //Wire declarations for instance 'op_8_54' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_54__in0;
  wire [15:0] op_8_54__in1;
  wire [15:0] op_8_54__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_54(
    .in0(op_8_54__in0),
    .in1(op_8_54__in1),
    .out(op_8_54__out)
  );

  //Wire declarations for instance 'op_8_55' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_55__in0;
  wire [15:0] op_8_55__in1;
  wire [15:0] op_8_55__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_55(
    .in0(op_8_55__in0),
    .in1(op_8_55__in1),
    .out(op_8_55__out)
  );

  //Wire declarations for instance 'op_8_56' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_56__in0;
  wire [15:0] op_8_56__in1;
  wire [15:0] op_8_56__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_56(
    .in0(op_8_56__in0),
    .in1(op_8_56__in1),
    .out(op_8_56__out)
  );

  //Wire declarations for instance 'op_8_57' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_57__in0;
  wire [15:0] op_8_57__in1;
  wire [15:0] op_8_57__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_57(
    .in0(op_8_57__in0),
    .in1(op_8_57__in1),
    .out(op_8_57__out)
  );

  //Wire declarations for instance 'op_8_58' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_58__in0;
  wire [15:0] op_8_58__in1;
  wire [15:0] op_8_58__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_58(
    .in0(op_8_58__in0),
    .in1(op_8_58__in1),
    .out(op_8_58__out)
  );

  //Wire declarations for instance 'op_8_59' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_59__in0;
  wire [15:0] op_8_59__in1;
  wire [15:0] op_8_59__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_59(
    .in0(op_8_59__in0),
    .in1(op_8_59__in1),
    .out(op_8_59__out)
  );

  //Wire declarations for instance 'op_8_6' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_6__in0;
  wire [15:0] op_8_6__in1;
  wire [15:0] op_8_6__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_6(
    .in0(op_8_6__in0),
    .in1(op_8_6__in1),
    .out(op_8_6__out)
  );

  //Wire declarations for instance 'op_8_60' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_60__in0;
  wire [15:0] op_8_60__in1;
  wire [15:0] op_8_60__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_60(
    .in0(op_8_60__in0),
    .in1(op_8_60__in1),
    .out(op_8_60__out)
  );

  //Wire declarations for instance 'op_8_61' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_61__in0;
  wire [15:0] op_8_61__in1;
  wire [15:0] op_8_61__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_61(
    .in0(op_8_61__in0),
    .in1(op_8_61__in1),
    .out(op_8_61__out)
  );

  //Wire declarations for instance 'op_8_62' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_62__in0;
  wire [15:0] op_8_62__in1;
  wire [15:0] op_8_62__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_62(
    .in0(op_8_62__in0),
    .in1(op_8_62__in1),
    .out(op_8_62__out)
  );

  //Wire declarations for instance 'op_8_63' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_63__in0;
  wire [15:0] op_8_63__in1;
  wire [15:0] op_8_63__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_63(
    .in0(op_8_63__in0),
    .in1(op_8_63__in1),
    .out(op_8_63__out)
  );

  //Wire declarations for instance 'op_8_64' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_64__in0;
  wire [15:0] op_8_64__in1;
  wire [15:0] op_8_64__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_64(
    .in0(op_8_64__in0),
    .in1(op_8_64__in1),
    .out(op_8_64__out)
  );

  //Wire declarations for instance 'op_8_65' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_65__in0;
  wire [15:0] op_8_65__in1;
  wire [15:0] op_8_65__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_65(
    .in0(op_8_65__in0),
    .in1(op_8_65__in1),
    .out(op_8_65__out)
  );

  //Wire declarations for instance 'op_8_66' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_66__in0;
  wire [15:0] op_8_66__in1;
  wire [15:0] op_8_66__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_66(
    .in0(op_8_66__in0),
    .in1(op_8_66__in1),
    .out(op_8_66__out)
  );

  //Wire declarations for instance 'op_8_67' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_67__in0;
  wire [15:0] op_8_67__in1;
  wire [15:0] op_8_67__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_67(
    .in0(op_8_67__in0),
    .in1(op_8_67__in1),
    .out(op_8_67__out)
  );

  //Wire declarations for instance 'op_8_68' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_68__in0;
  wire [15:0] op_8_68__in1;
  wire [15:0] op_8_68__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_68(
    .in0(op_8_68__in0),
    .in1(op_8_68__in1),
    .out(op_8_68__out)
  );

  //Wire declarations for instance 'op_8_69' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_69__in0;
  wire [15:0] op_8_69__in1;
  wire [15:0] op_8_69__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_69(
    .in0(op_8_69__in0),
    .in1(op_8_69__in1),
    .out(op_8_69__out)
  );

  //Wire declarations for instance 'op_8_7' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_7__in0;
  wire [15:0] op_8_7__in1;
  wire [15:0] op_8_7__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_7(
    .in0(op_8_7__in0),
    .in1(op_8_7__in1),
    .out(op_8_7__out)
  );

  //Wire declarations for instance 'op_8_70' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_70__in0;
  wire [15:0] op_8_70__in1;
  wire [15:0] op_8_70__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_70(
    .in0(op_8_70__in0),
    .in1(op_8_70__in1),
    .out(op_8_70__out)
  );

  //Wire declarations for instance 'op_8_71' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_71__in0;
  wire [15:0] op_8_71__in1;
  wire [15:0] op_8_71__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_71(
    .in0(op_8_71__in0),
    .in1(op_8_71__in1),
    .out(op_8_71__out)
  );

  //Wire declarations for instance 'op_8_72' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_72__in0;
  wire [15:0] op_8_72__in1;
  wire [15:0] op_8_72__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_72(
    .in0(op_8_72__in0),
    .in1(op_8_72__in1),
    .out(op_8_72__out)
  );

  //Wire declarations for instance 'op_8_73' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_73__in0;
  wire [15:0] op_8_73__in1;
  wire [15:0] op_8_73__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_73(
    .in0(op_8_73__in0),
    .in1(op_8_73__in1),
    .out(op_8_73__out)
  );

  //Wire declarations for instance 'op_8_74' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_74__in0;
  wire [15:0] op_8_74__in1;
  wire [15:0] op_8_74__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_74(
    .in0(op_8_74__in0),
    .in1(op_8_74__in1),
    .out(op_8_74__out)
  );

  //Wire declarations for instance 'op_8_75' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_75__in0;
  wire [15:0] op_8_75__in1;
  wire [15:0] op_8_75__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_75(
    .in0(op_8_75__in0),
    .in1(op_8_75__in1),
    .out(op_8_75__out)
  );

  //Wire declarations for instance 'op_8_76' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_76__in0;
  wire [15:0] op_8_76__in1;
  wire [15:0] op_8_76__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_76(
    .in0(op_8_76__in0),
    .in1(op_8_76__in1),
    .out(op_8_76__out)
  );

  //Wire declarations for instance 'op_8_77' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_77__in0;
  wire [15:0] op_8_77__in1;
  wire [15:0] op_8_77__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_77(
    .in0(op_8_77__in0),
    .in1(op_8_77__in1),
    .out(op_8_77__out)
  );

  //Wire declarations for instance 'op_8_78' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_78__in0;
  wire [15:0] op_8_78__in1;
  wire [15:0] op_8_78__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_78(
    .in0(op_8_78__in0),
    .in1(op_8_78__in1),
    .out(op_8_78__out)
  );

  //Wire declarations for instance 'op_8_79' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_79__in0;
  wire [15:0] op_8_79__in1;
  wire [15:0] op_8_79__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_79(
    .in0(op_8_79__in0),
    .in1(op_8_79__in1),
    .out(op_8_79__out)
  );

  //Wire declarations for instance 'op_8_8' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_8__in0;
  wire [15:0] op_8_8__in1;
  wire [15:0] op_8_8__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_8(
    .in0(op_8_8__in0),
    .in1(op_8_8__in1),
    .out(op_8_8__out)
  );

  //Wire declarations for instance 'op_8_80' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_80__in0;
  wire [15:0] op_8_80__in1;
  wire [15:0] op_8_80__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_80(
    .in0(op_8_80__in0),
    .in1(op_8_80__in1),
    .out(op_8_80__out)
  );

  //Wire declarations for instance 'op_8_81' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_81__in0;
  wire [15:0] op_8_81__in1;
  wire [15:0] op_8_81__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_81(
    .in0(op_8_81__in0),
    .in1(op_8_81__in1),
    .out(op_8_81__out)
  );

  //Wire declarations for instance 'op_8_82' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_82__in0;
  wire [15:0] op_8_82__in1;
  wire [15:0] op_8_82__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_82(
    .in0(op_8_82__in0),
    .in1(op_8_82__in1),
    .out(op_8_82__out)
  );

  //Wire declarations for instance 'op_8_83' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_83__in0;
  wire [15:0] op_8_83__in1;
  wire [15:0] op_8_83__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_83(
    .in0(op_8_83__in0),
    .in1(op_8_83__in1),
    .out(op_8_83__out)
  );

  //Wire declarations for instance 'op_8_84' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_84__in0;
  wire [15:0] op_8_84__in1;
  wire [15:0] op_8_84__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_84(
    .in0(op_8_84__in0),
    .in1(op_8_84__in1),
    .out(op_8_84__out)
  );

  //Wire declarations for instance 'op_8_85' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_85__in0;
  wire [15:0] op_8_85__in1;
  wire [15:0] op_8_85__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_85(
    .in0(op_8_85__in0),
    .in1(op_8_85__in1),
    .out(op_8_85__out)
  );

  //Wire declarations for instance 'op_8_86' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_86__in0;
  wire [15:0] op_8_86__in1;
  wire [15:0] op_8_86__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_86(
    .in0(op_8_86__in0),
    .in1(op_8_86__in1),
    .out(op_8_86__out)
  );

  //Wire declarations for instance 'op_8_87' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_87__in0;
  wire [15:0] op_8_87__in1;
  wire [15:0] op_8_87__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_87(
    .in0(op_8_87__in0),
    .in1(op_8_87__in1),
    .out(op_8_87__out)
  );

  //Wire declarations for instance 'op_8_88' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_88__in0;
  wire [15:0] op_8_88__in1;
  wire [15:0] op_8_88__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_88(
    .in0(op_8_88__in0),
    .in1(op_8_88__in1),
    .out(op_8_88__out)
  );

  //Wire declarations for instance 'op_8_89' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_89__in0;
  wire [15:0] op_8_89__in1;
  wire [15:0] op_8_89__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_89(
    .in0(op_8_89__in0),
    .in1(op_8_89__in1),
    .out(op_8_89__out)
  );

  //Wire declarations for instance 'op_8_9' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_9__in0;
  wire [15:0] op_8_9__in1;
  wire [15:0] op_8_9__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_9(
    .in0(op_8_9__in0),
    .in1(op_8_9__in1),
    .out(op_8_9__out)
  );

  //Wire declarations for instance 'op_8_90' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_90__in0;
  wire [15:0] op_8_90__in1;
  wire [15:0] op_8_90__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_90(
    .in0(op_8_90__in0),
    .in1(op_8_90__in1),
    .out(op_8_90__out)
  );

  //Wire declarations for instance 'op_8_91' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_91__in0;
  wire [15:0] op_8_91__in1;
  wire [15:0] op_8_91__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_91(
    .in0(op_8_91__in0),
    .in1(op_8_91__in1),
    .out(op_8_91__out)
  );

  //Wire declarations for instance 'op_8_92' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_92__in0;
  wire [15:0] op_8_92__in1;
  wire [15:0] op_8_92__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_92(
    .in0(op_8_92__in0),
    .in1(op_8_92__in1),
    .out(op_8_92__out)
  );

  //Wire declarations for instance 'op_8_93' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_93__in0;
  wire [15:0] op_8_93__in1;
  wire [15:0] op_8_93__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_93(
    .in0(op_8_93__in0),
    .in1(op_8_93__in1),
    .out(op_8_93__out)
  );

  //Wire declarations for instance 'op_8_94' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_94__in0;
  wire [15:0] op_8_94__in1;
  wire [15:0] op_8_94__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_94(
    .in0(op_8_94__in0),
    .in1(op_8_94__in1),
    .out(op_8_94__out)
  );

  //Wire declarations for instance 'op_8_95' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_95__in0;
  wire [15:0] op_8_95__in1;
  wire [15:0] op_8_95__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_95(
    .in0(op_8_95__in0),
    .in1(op_8_95__in1),
    .out(op_8_95__out)
  );

  //Wire declarations for instance 'op_8_96' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_96__in0;
  wire [15:0] op_8_96__in1;
  wire [15:0] op_8_96__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_96(
    .in0(op_8_96__in0),
    .in1(op_8_96__in1),
    .out(op_8_96__out)
  );

  //Wire declarations for instance 'op_8_97' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_97__in0;
  wire [15:0] op_8_97__in1;
  wire [15:0] op_8_97__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_97(
    .in0(op_8_97__in0),
    .in1(op_8_97__in1),
    .out(op_8_97__out)
  );

  //Wire declarations for instance 'op_8_98' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_98__in0;
  wire [15:0] op_8_98__in1;
  wire [15:0] op_8_98__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_98(
    .in0(op_8_98__in0),
    .in1(op_8_98__in1),
    .out(op_8_98__out)
  );

  //Wire declarations for instance 'op_8_99' (Module renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___)
  wire [15:0] op_8_99__in0;
  wire [15:0] op_8_99__in1;
  wire [15:0] op_8_99__out;
  renamedForReduce_opAdd16_I0_In_Bits_16___I1_In_Bits_16___O_Out_Bits_16___ op_8_99(
    .in0(op_8_99__in0),
    .in1(op_8_99__in1),
    .out(op_8_99__out)
  );

  //All the connections
  assign out[15:0] = op_0_0__out[15:0];
  assign op_0_0__in0[15:0] = op_1_0__out[15:0];
  assign op_0_0__in1[15:0] = op_1_1__out[15:0];
  assign op_1_0__in0[15:0] = op_2_0__out[15:0];
  assign op_1_0__in1[15:0] = op_2_1__out[15:0];
  assign op_1_1__in0[15:0] = op_2_2__out[15:0];
  assign op_1_1__in1[15:0] = op_2_3__out[15:0];
  assign op_2_0__in0[15:0] = op_3_0__out[15:0];
  assign op_2_0__in1[15:0] = op_3_1__out[15:0];
  assign op_2_1__in0[15:0] = op_3_2__out[15:0];
  assign op_2_1__in1[15:0] = op_3_3__out[15:0];
  assign op_2_2__in0[15:0] = op_3_4__out[15:0];
  assign op_2_2__in1[15:0] = op_3_5__out[15:0];
  assign op_2_3__in0[15:0] = op_3_6__out[15:0];
  assign op_2_3__in1[15:0] = op_3_7__out[15:0];
  assign op_3_0__in0[15:0] = op_4_0__out[15:0];
  assign op_3_0__in1[15:0] = op_4_1__out[15:0];
  assign op_3_1__in0[15:0] = op_4_2__out[15:0];
  assign op_3_1__in1[15:0] = op_4_3__out[15:0];
  assign op_3_2__in0[15:0] = op_4_4__out[15:0];
  assign op_3_2__in1[15:0] = op_4_5__out[15:0];
  assign op_3_3__in0[15:0] = op_4_6__out[15:0];
  assign op_3_3__in1[15:0] = op_4_7__out[15:0];
  assign op_3_4__in0[15:0] = op_4_8__out[15:0];
  assign op_3_4__in1[15:0] = op_4_9__out[15:0];
  assign op_3_5__in0[15:0] = op_4_10__out[15:0];
  assign op_3_5__in1[15:0] = op_4_11__out[15:0];
  assign op_3_6__in0[15:0] = op_4_12__out[15:0];
  assign op_3_6__in1[15:0] = op_4_13__out[15:0];
  assign op_3_7__in0[15:0] = op_4_14__out[15:0];
  assign op_3_7__in1[15:0] = op_4_15__out[15:0];
  assign op_4_0__in0[15:0] = op_5_0__out[15:0];
  assign op_4_0__in1[15:0] = op_5_1__out[15:0];
  assign op_4_1__in0[15:0] = op_5_2__out[15:0];
  assign op_4_1__in1[15:0] = op_5_3__out[15:0];
  assign op_4_2__in0[15:0] = op_5_4__out[15:0];
  assign op_4_2__in1[15:0] = op_5_5__out[15:0];
  assign op_4_3__in0[15:0] = op_5_6__out[15:0];
  assign op_4_3__in1[15:0] = op_5_7__out[15:0];
  assign op_4_4__in0[15:0] = op_5_8__out[15:0];
  assign op_4_4__in1[15:0] = op_5_9__out[15:0];
  assign op_4_5__in0[15:0] = op_5_10__out[15:0];
  assign op_4_5__in1[15:0] = op_5_11__out[15:0];
  assign op_4_6__in0[15:0] = op_5_12__out[15:0];
  assign op_4_6__in1[15:0] = op_5_13__out[15:0];
  assign op_4_7__in0[15:0] = op_5_14__out[15:0];
  assign op_5_16__in1[15:0] = op_6_33__out[15:0];
  assign op_4_7__in1[15:0] = op_5_15__out[15:0];
  assign op_4_8__in0[15:0] = op_5_16__out[15:0];
  assign op_4_8__in1[15:0] = op_5_17__out[15:0];
  assign op_4_9__in0[15:0] = op_5_18__out[15:0];
  assign op_4_9__in1[15:0] = op_5_19__out[15:0];
  assign op_4_10__in0[15:0] = op_5_20__out[15:0];
  assign op_4_10__in1[15:0] = op_5_21__out[15:0];
  assign op_4_11__in0[15:0] = op_5_22__out[15:0];
  assign op_4_11__in1[15:0] = op_5_23__out[15:0];
  assign op_4_12__in0[15:0] = op_5_24__out[15:0];
  assign op_4_12__in1[15:0] = op_5_25__out[15:0];
  assign op_4_13__in0[15:0] = op_5_26__out[15:0];
  assign op_4_13__in1[15:0] = op_5_27__out[15:0];
  assign op_4_14__in0[15:0] = op_5_28__out[15:0];
  assign op_4_14__in1[15:0] = op_5_29__out[15:0];
  assign op_4_15__in0[15:0] = op_5_30__out[15:0];
  assign op_4_15__in1[15:0] = op_5_31__out[15:0];
  assign op_5_0__in0[15:0] = op_6_0__out[15:0];
  assign op_5_0__in1[15:0] = op_6_1__out[15:0];
  assign op_5_1__in0[15:0] = op_6_2__out[15:0];
  assign op_5_1__in1[15:0] = op_6_3__out[15:0];
  assign op_5_2__in0[15:0] = op_6_4__out[15:0];
  assign op_5_2__in1[15:0] = op_6_5__out[15:0];
  assign op_5_3__in0[15:0] = op_6_6__out[15:0];
  assign op_5_3__in1[15:0] = op_6_7__out[15:0];
  assign op_5_4__in0[15:0] = op_6_8__out[15:0];
  assign op_5_4__in1[15:0] = op_6_9__out[15:0];
  assign op_5_5__in0[15:0] = op_6_10__out[15:0];
  assign op_5_5__in1[15:0] = op_6_11__out[15:0];
  assign op_5_6__in0[15:0] = op_6_12__out[15:0];
  assign op_5_6__in1[15:0] = op_6_13__out[15:0];
  assign op_5_7__in0[15:0] = op_6_14__out[15:0];
  assign op_5_7__in1[15:0] = op_6_15__out[15:0];
  assign op_5_8__in0[15:0] = op_6_16__out[15:0];
  assign op_5_8__in1[15:0] = op_6_17__out[15:0];
  assign op_5_9__in0[15:0] = op_6_18__out[15:0];
  assign op_5_9__in1[15:0] = op_6_19__out[15:0];
  assign op_5_10__in0[15:0] = op_6_20__out[15:0];
  assign op_5_10__in1[15:0] = op_6_21__out[15:0];
  assign op_5_11__in0[15:0] = op_6_22__out[15:0];
  assign op_5_11__in1[15:0] = op_6_23__out[15:0];
  assign op_5_12__in0[15:0] = op_6_24__out[15:0];
  assign op_5_12__in1[15:0] = op_6_25__out[15:0];
  assign op_5_13__in0[15:0] = op_6_26__out[15:0];
  assign op_5_13__in1[15:0] = op_6_27__out[15:0];
  assign op_5_14__in0[15:0] = op_6_28__out[15:0];
  assign op_5_14__in1[15:0] = op_6_29__out[15:0];
  assign op_5_15__in0[15:0] = op_6_30__out[15:0];
  assign op_5_15__in1[15:0] = op_6_31__out[15:0];
  assign op_5_16__in0[15:0] = op_6_32__out[15:0];
  assign op_6_35__in1[15:0] = op_7_71__out[15:0];
  assign op_5_17__in0[15:0] = op_6_34__out[15:0];
  assign op_5_17__in1[15:0] = op_6_35__out[15:0];
  assign op_5_18__in0[15:0] = op_6_36__out[15:0];
  assign op_5_18__in1[15:0] = op_6_37__out[15:0];
  assign op_5_19__in0[15:0] = op_6_38__out[15:0];
  assign op_5_19__in1[15:0] = op_6_39__out[15:0];
  assign op_5_20__in0[15:0] = op_6_40__out[15:0];
  assign op_5_20__in1[15:0] = op_6_41__out[15:0];
  assign op_5_21__in0[15:0] = op_6_42__out[15:0];
  assign op_5_21__in1[15:0] = op_6_43__out[15:0];
  assign op_5_22__in0[15:0] = op_6_44__out[15:0];
  assign op_5_22__in1[15:0] = op_6_45__out[15:0];
  assign op_5_23__in0[15:0] = op_6_46__out[15:0];
  assign op_5_23__in1[15:0] = op_6_47__out[15:0];
  assign op_5_24__in0[15:0] = op_6_48__out[15:0];
  assign op_5_24__in1[15:0] = op_6_49__out[15:0];
  assign op_5_25__in0[15:0] = op_6_50__out[15:0];
  assign op_5_25__in1[15:0] = op_6_51__out[15:0];
  assign op_5_26__in0[15:0] = op_6_52__out[15:0];
  assign op_5_26__in1[15:0] = op_6_53__out[15:0];
  assign op_5_27__in0[15:0] = op_6_54__out[15:0];
  assign op_5_27__in1[15:0] = op_6_55__out[15:0];
  assign op_5_28__in0[15:0] = op_6_56__out[15:0];
  assign op_5_28__in1[15:0] = op_6_57__out[15:0];
  assign op_5_29__in0[15:0] = op_6_58__out[15:0];
  assign op_5_29__in1[15:0] = op_6_59__out[15:0];
  assign op_5_30__in0[15:0] = op_6_60__out[15:0];
  assign op_5_30__in1[15:0] = op_6_61__out[15:0];
  assign op_5_31__in0[15:0] = op_6_62__out[15:0];
  assign op_5_31__in1[15:0] = op_6_63__out[15:0];
  assign op_6_0__in0[15:0] = op_7_0__out[15:0];
  assign op_6_0__in1[15:0] = op_7_1__out[15:0];
  assign op_6_1__in0[15:0] = op_7_2__out[15:0];
  assign op_6_1__in1[15:0] = op_7_3__out[15:0];
  assign op_6_2__in0[15:0] = op_7_4__out[15:0];
  assign op_6_2__in1[15:0] = op_7_5__out[15:0];
  assign op_6_3__in0[15:0] = op_7_6__out[15:0];
  assign op_6_3__in1[15:0] = op_7_7__out[15:0];
  assign op_6_4__in0[15:0] = op_7_8__out[15:0];
  assign op_6_4__in1[15:0] = op_7_9__out[15:0];
  assign op_6_5__in0[15:0] = op_7_10__out[15:0];
  assign op_6_5__in1[15:0] = op_7_11__out[15:0];
  assign op_6_6__in0[15:0] = op_7_12__out[15:0];
  assign op_6_6__in1[15:0] = op_7_13__out[15:0];
  assign op_6_7__in0[15:0] = op_7_14__out[15:0];
  assign op_6_7__in1[15:0] = op_7_15__out[15:0];
  assign op_6_8__in0[15:0] = op_7_16__out[15:0];
  assign op_6_8__in1[15:0] = op_7_17__out[15:0];
  assign op_6_9__in0[15:0] = op_7_18__out[15:0];
  assign op_6_9__in1[15:0] = op_7_19__out[15:0];
  assign op_6_10__in0[15:0] = op_7_20__out[15:0];
  assign op_6_10__in1[15:0] = op_7_21__out[15:0];
  assign op_6_11__in0[15:0] = op_7_22__out[15:0];
  assign op_6_11__in1[15:0] = op_7_23__out[15:0];
  assign op_6_12__in0[15:0] = op_7_24__out[15:0];
  assign op_6_12__in1[15:0] = op_7_25__out[15:0];
  assign op_6_13__in0[15:0] = op_7_26__out[15:0];
  assign op_6_13__in1[15:0] = op_7_27__out[15:0];
  assign op_6_14__in0[15:0] = op_7_28__out[15:0];
  assign op_6_14__in1[15:0] = op_7_29__out[15:0];
  assign op_6_15__in0[15:0] = op_7_30__out[15:0];
  assign op_6_15__in1[15:0] = op_7_31__out[15:0];
  assign op_6_16__in0[15:0] = op_7_32__out[15:0];
  assign op_6_16__in1[15:0] = op_7_33__out[15:0];
  assign op_6_17__in0[15:0] = op_7_34__out[15:0];
  assign op_6_17__in1[15:0] = op_7_35__out[15:0];
  assign op_6_18__in0[15:0] = op_7_36__out[15:0];
  assign op_6_18__in1[15:0] = op_7_37__out[15:0];
  assign op_6_19__in0[15:0] = op_7_38__out[15:0];
  assign op_6_19__in1[15:0] = op_7_39__out[15:0];
  assign op_6_20__in0[15:0] = op_7_40__out[15:0];
  assign op_6_20__in1[15:0] = op_7_41__out[15:0];
  assign op_6_21__in0[15:0] = op_7_42__out[15:0];
  assign op_6_21__in1[15:0] = op_7_43__out[15:0];
  assign op_6_22__in0[15:0] = op_7_44__out[15:0];
  assign op_6_22__in1[15:0] = op_7_45__out[15:0];
  assign op_6_23__in0[15:0] = op_7_46__out[15:0];
  assign op_6_23__in1[15:0] = op_7_47__out[15:0];
  assign op_6_24__in0[15:0] = op_7_48__out[15:0];
  assign op_6_24__in1[15:0] = op_7_49__out[15:0];
  assign op_6_25__in0[15:0] = op_7_50__out[15:0];
  assign op_6_25__in1[15:0] = op_7_51__out[15:0];
  assign op_6_26__in0[15:0] = op_7_52__out[15:0];
  assign op_6_26__in1[15:0] = op_7_53__out[15:0];
  assign op_6_27__in0[15:0] = op_7_54__out[15:0];
  assign op_6_27__in1[15:0] = op_7_55__out[15:0];
  assign op_6_28__in0[15:0] = op_7_56__out[15:0];
  assign op_6_28__in1[15:0] = op_7_57__out[15:0];
  assign op_6_29__in0[15:0] = op_7_58__out[15:0];
  assign op_6_29__in1[15:0] = op_7_59__out[15:0];
  assign op_6_30__in0[15:0] = op_7_60__out[15:0];
  assign op_6_30__in1[15:0] = op_7_61__out[15:0];
  assign op_6_31__in0[15:0] = op_7_62__out[15:0];
  assign op_6_31__in1[15:0] = op_7_63__out[15:0];
  assign op_6_32__in0[15:0] = op_7_64__out[15:0];
  assign op_6_32__in1[15:0] = op_7_65__out[15:0];
  assign op_6_33__in0[15:0] = op_7_66__out[15:0];
  assign op_6_33__in1[15:0] = op_7_67__out[15:0];
  assign op_6_34__in0[15:0] = op_7_68__out[15:0];
  assign op_6_34__in1[15:0] = op_7_69__out[15:0];
  assign op_6_35__in0[15:0] = op_7_70__out[15:0];
  assign op_8_153__in0[15:0] = in_306[15:0];
  assign op_7_76__in1[15:0] = op_8_153__out[15:0];
  assign op_8_153__in1[15:0] = in_307[15:0];
  assign op_6_36__in0[15:0] = op_7_72__out[15:0];
  assign op_6_36__in1[15:0] = op_7_73__out[15:0];
  assign op_6_37__in0[15:0] = op_7_74__out[15:0];
  assign op_6_37__in1[15:0] = op_7_75__out[15:0];
  assign op_6_38__in0[15:0] = op_7_76__out[15:0];
  assign op_6_38__in1[15:0] = op_7_77__out[15:0];
  assign op_6_39__in0[15:0] = op_7_78__out[15:0];
  assign op_6_39__in1[15:0] = op_7_79__out[15:0];
  assign op_6_40__in0[15:0] = op_7_80__out[15:0];
  assign op_6_40__in1[15:0] = op_7_81__out[15:0];
  assign op_6_41__in0[15:0] = op_7_82__out[15:0];
  assign op_6_41__in1[15:0] = op_7_83__out[15:0];
  assign op_6_42__in0[15:0] = op_7_84__out[15:0];
  assign op_6_42__in1[15:0] = op_7_85__out[15:0];
  assign op_6_43__in0[15:0] = op_7_86__out[15:0];
  assign op_6_43__in1[15:0] = op_7_87__out[15:0];
  assign op_6_44__in0[15:0] = op_7_88__out[15:0];
  assign op_6_44__in1[15:0] = op_7_89__out[15:0];
  assign op_6_45__in0[15:0] = op_7_90__out[15:0];
  assign op_6_45__in1[15:0] = op_7_91__out[15:0];
  assign op_6_46__in0[15:0] = op_7_92__out[15:0];
  assign op_6_46__in1[15:0] = op_7_93__out[15:0];
  assign op_6_47__in0[15:0] = op_7_94__out[15:0];
  assign op_6_47__in1[15:0] = op_7_95__out[15:0];
  assign op_6_48__in0[15:0] = op_7_96__out[15:0];
  assign op_6_48__in1[15:0] = op_7_97__out[15:0];
  assign op_6_49__in0[15:0] = op_7_98__out[15:0];
  assign op_6_49__in1[15:0] = op_7_99__out[15:0];
  assign op_6_50__in0[15:0] = op_7_100__out[15:0];
  assign op_6_50__in1[15:0] = op_7_101__out[15:0];
  assign op_6_51__in0[15:0] = op_7_102__out[15:0];
  assign op_6_51__in1[15:0] = op_7_103__out[15:0];
  assign op_6_52__in0[15:0] = op_7_104__out[15:0];
  assign op_6_52__in1[15:0] = op_7_105__out[15:0];
  assign op_6_53__in0[15:0] = op_7_106__out[15:0];
  assign op_6_53__in1[15:0] = op_7_107__out[15:0];
  assign op_6_54__in0[15:0] = op_7_108__out[15:0];
  assign op_6_54__in1[15:0] = op_7_109__out[15:0];
  assign op_6_55__in0[15:0] = op_7_110__out[15:0];
  assign op_6_55__in1[15:0] = op_7_111__out[15:0];
  assign op_6_56__in0[15:0] = op_7_112__out[15:0];
  assign op_6_56__in1[15:0] = op_7_113__out[15:0];
  assign op_6_57__in0[15:0] = op_7_114__out[15:0];
  assign op_6_57__in1[15:0] = op_7_115__out[15:0];
  assign op_6_58__in0[15:0] = op_7_116__out[15:0];
  assign op_6_58__in1[15:0] = op_7_117__out[15:0];
  assign op_6_59__in0[15:0] = op_7_118__out[15:0];
  assign op_6_59__in1[15:0] = op_7_119__out[15:0];
  assign op_6_60__in0[15:0] = op_7_120__out[15:0];
  assign op_6_60__in1[15:0] = op_7_121__out[15:0];
  assign op_6_61__in0[15:0] = op_7_122__out[15:0];
  assign op_6_61__in1[15:0] = op_7_123__out[15:0];
  assign op_6_62__in0[15:0] = op_7_124__out[15:0];
  assign op_6_62__in1[15:0] = op_7_125__out[15:0];
  assign op_6_63__in0[15:0] = op_7_126__out[15:0];
  assign op_6_63__in1[15:0] = op_7_127__out[15:0];
  assign op_8_0__in1[15:0] = in_1[15:0];
  assign op_8_0__in0[15:0] = in_0[15:0];
  assign op_7_0__in0[15:0] = op_8_0__out[15:0];
  assign op_8_1__in1[15:0] = in_3[15:0];
  assign op_8_1__in0[15:0] = in_2[15:0];
  assign op_7_0__in1[15:0] = op_8_1__out[15:0];
  assign op_8_2__in1[15:0] = in_5[15:0];
  assign op_8_2__in0[15:0] = in_4[15:0];
  assign op_7_1__in0[15:0] = op_8_2__out[15:0];
  assign op_8_3__in1[15:0] = in_7[15:0];
  assign op_8_3__in0[15:0] = in_6[15:0];
  assign op_7_1__in1[15:0] = op_8_3__out[15:0];
  assign op_8_4__in1[15:0] = in_9[15:0];
  assign op_8_4__in0[15:0] = in_8[15:0];
  assign op_7_2__in0[15:0] = op_8_4__out[15:0];
  assign op_8_5__in1[15:0] = in_11[15:0];
  assign op_8_5__in0[15:0] = in_10[15:0];
  assign op_7_2__in1[15:0] = op_8_5__out[15:0];
  assign op_8_6__in1[15:0] = in_13[15:0];
  assign op_8_6__in0[15:0] = in_12[15:0];
  assign op_7_3__in0[15:0] = op_8_6__out[15:0];
  assign op_8_7__in1[15:0] = in_15[15:0];
  assign op_8_7__in0[15:0] = in_14[15:0];
  assign op_7_3__in1[15:0] = op_8_7__out[15:0];
  assign op_8_8__in1[15:0] = in_17[15:0];
  assign op_8_8__in0[15:0] = in_16[15:0];
  assign op_7_4__in0[15:0] = op_8_8__out[15:0];
  assign op_8_9__in1[15:0] = in_19[15:0];
  assign op_8_9__in0[15:0] = in_18[15:0];
  assign op_7_4__in1[15:0] = op_8_9__out[15:0];
  assign op_8_10__in1[15:0] = in_21[15:0];
  assign op_8_10__in0[15:0] = in_20[15:0];
  assign op_7_5__in0[15:0] = op_8_10__out[15:0];
  assign op_8_11__in1[15:0] = in_23[15:0];
  assign op_8_11__in0[15:0] = in_22[15:0];
  assign op_7_5__in1[15:0] = op_8_11__out[15:0];
  assign op_8_12__in1[15:0] = in_25[15:0];
  assign op_8_12__in0[15:0] = in_24[15:0];
  assign op_7_6__in0[15:0] = op_8_12__out[15:0];
  assign op_8_13__in1[15:0] = in_27[15:0];
  assign op_8_13__in0[15:0] = in_26[15:0];
  assign op_7_6__in1[15:0] = op_8_13__out[15:0];
  assign op_8_14__in1[15:0] = in_29[15:0];
  assign op_8_14__in0[15:0] = in_28[15:0];
  assign op_7_7__in0[15:0] = op_8_14__out[15:0];
  assign op_8_15__in1[15:0] = in_31[15:0];
  assign op_8_15__in0[15:0] = in_30[15:0];
  assign op_7_7__in1[15:0] = op_8_15__out[15:0];
  assign op_8_16__in1[15:0] = in_33[15:0];
  assign op_8_16__in0[15:0] = in_32[15:0];
  assign op_7_8__in0[15:0] = op_8_16__out[15:0];
  assign op_8_17__in1[15:0] = in_35[15:0];
  assign op_8_17__in0[15:0] = in_34[15:0];
  assign op_7_8__in1[15:0] = op_8_17__out[15:0];
  assign op_8_18__in1[15:0] = in_37[15:0];
  assign op_8_18__in0[15:0] = in_36[15:0];
  assign op_7_9__in0[15:0] = op_8_18__out[15:0];
  assign op_8_19__in1[15:0] = in_39[15:0];
  assign op_8_19__in0[15:0] = in_38[15:0];
  assign op_7_9__in1[15:0] = op_8_19__out[15:0];
  assign op_8_20__in1[15:0] = in_41[15:0];
  assign op_8_20__in0[15:0] = in_40[15:0];
  assign op_7_10__in0[15:0] = op_8_20__out[15:0];
  assign op_8_21__in1[15:0] = in_43[15:0];
  assign op_8_21__in0[15:0] = in_42[15:0];
  assign op_7_10__in1[15:0] = op_8_21__out[15:0];
  assign op_8_22__in1[15:0] = in_45[15:0];
  assign op_8_22__in0[15:0] = in_44[15:0];
  assign op_7_11__in0[15:0] = op_8_22__out[15:0];
  assign op_8_23__in1[15:0] = in_47[15:0];
  assign op_8_23__in0[15:0] = in_46[15:0];
  assign op_7_11__in1[15:0] = op_8_23__out[15:0];
  assign op_8_24__in1[15:0] = in_49[15:0];
  assign op_8_24__in0[15:0] = in_48[15:0];
  assign op_7_12__in0[15:0] = op_8_24__out[15:0];
  assign op_8_25__in1[15:0] = in_51[15:0];
  assign op_8_25__in0[15:0] = in_50[15:0];
  assign op_7_12__in1[15:0] = op_8_25__out[15:0];
  assign op_8_26__in1[15:0] = in_53[15:0];
  assign op_8_26__in0[15:0] = in_52[15:0];
  assign op_7_13__in0[15:0] = op_8_26__out[15:0];
  assign op_8_27__in1[15:0] = in_55[15:0];
  assign op_8_27__in0[15:0] = in_54[15:0];
  assign op_7_13__in1[15:0] = op_8_27__out[15:0];
  assign op_8_28__in1[15:0] = in_57[15:0];
  assign op_8_28__in0[15:0] = in_56[15:0];
  assign op_7_14__in0[15:0] = op_8_28__out[15:0];
  assign op_8_29__in1[15:0] = in_59[15:0];
  assign op_8_29__in0[15:0] = in_58[15:0];
  assign op_7_14__in1[15:0] = op_8_29__out[15:0];
  assign op_8_30__in1[15:0] = in_61[15:0];
  assign op_8_30__in0[15:0] = in_60[15:0];
  assign op_7_15__in0[15:0] = op_8_30__out[15:0];
  assign op_8_31__in1[15:0] = in_63[15:0];
  assign op_8_31__in0[15:0] = in_62[15:0];
  assign op_7_15__in1[15:0] = op_8_31__out[15:0];
  assign op_8_32__in1[15:0] = in_65[15:0];
  assign op_8_32__in0[15:0] = in_64[15:0];
  assign op_7_16__in0[15:0] = op_8_32__out[15:0];
  assign op_8_33__in1[15:0] = in_67[15:0];
  assign op_8_33__in0[15:0] = in_66[15:0];
  assign op_7_16__in1[15:0] = op_8_33__out[15:0];
  assign op_8_34__in1[15:0] = in_69[15:0];
  assign op_8_34__in0[15:0] = in_68[15:0];
  assign op_7_17__in0[15:0] = op_8_34__out[15:0];
  assign op_8_35__in1[15:0] = in_71[15:0];
  assign op_8_35__in0[15:0] = in_70[15:0];
  assign op_7_17__in1[15:0] = op_8_35__out[15:0];
  assign op_8_36__in1[15:0] = in_73[15:0];
  assign op_8_36__in0[15:0] = in_72[15:0];
  assign op_7_18__in0[15:0] = op_8_36__out[15:0];
  assign op_8_37__in1[15:0] = in_75[15:0];
  assign op_8_37__in0[15:0] = in_74[15:0];
  assign op_7_18__in1[15:0] = op_8_37__out[15:0];
  assign op_8_38__in1[15:0] = in_77[15:0];
  assign op_8_38__in0[15:0] = in_76[15:0];
  assign op_7_19__in0[15:0] = op_8_38__out[15:0];
  assign op_8_39__in1[15:0] = in_79[15:0];
  assign op_8_39__in0[15:0] = in_78[15:0];
  assign op_7_19__in1[15:0] = op_8_39__out[15:0];
  assign op_8_40__in1[15:0] = in_81[15:0];
  assign op_8_40__in0[15:0] = in_80[15:0];
  assign op_7_20__in0[15:0] = op_8_40__out[15:0];
  assign op_8_41__in1[15:0] = in_83[15:0];
  assign op_8_41__in0[15:0] = in_82[15:0];
  assign op_7_20__in1[15:0] = op_8_41__out[15:0];
  assign op_8_42__in1[15:0] = in_85[15:0];
  assign op_8_42__in0[15:0] = in_84[15:0];
  assign op_7_21__in0[15:0] = op_8_42__out[15:0];
  assign op_8_43__in1[15:0] = in_87[15:0];
  assign op_8_43__in0[15:0] = in_86[15:0];
  assign op_7_21__in1[15:0] = op_8_43__out[15:0];
  assign op_8_44__in1[15:0] = in_89[15:0];
  assign op_8_44__in0[15:0] = in_88[15:0];
  assign op_7_22__in0[15:0] = op_8_44__out[15:0];
  assign op_8_45__in1[15:0] = in_91[15:0];
  assign op_8_45__in0[15:0] = in_90[15:0];
  assign op_7_22__in1[15:0] = op_8_45__out[15:0];
  assign op_8_46__in1[15:0] = in_93[15:0];
  assign op_8_46__in0[15:0] = in_92[15:0];
  assign op_7_23__in0[15:0] = op_8_46__out[15:0];
  assign op_8_47__in1[15:0] = in_95[15:0];
  assign op_8_47__in0[15:0] = in_94[15:0];
  assign op_7_23__in1[15:0] = op_8_47__out[15:0];
  assign op_8_48__in1[15:0] = in_97[15:0];
  assign op_8_48__in0[15:0] = in_96[15:0];
  assign op_7_24__in0[15:0] = op_8_48__out[15:0];
  assign op_8_49__in1[15:0] = in_99[15:0];
  assign op_8_49__in0[15:0] = in_98[15:0];
  assign op_7_24__in1[15:0] = op_8_49__out[15:0];
  assign op_8_50__in1[15:0] = in_101[15:0];
  assign op_8_50__in0[15:0] = in_100[15:0];
  assign op_7_25__in0[15:0] = op_8_50__out[15:0];
  assign op_8_51__in1[15:0] = in_103[15:0];
  assign op_8_51__in0[15:0] = in_102[15:0];
  assign op_7_25__in1[15:0] = op_8_51__out[15:0];
  assign op_8_52__in1[15:0] = in_105[15:0];
  assign op_8_52__in0[15:0] = in_104[15:0];
  assign op_7_26__in0[15:0] = op_8_52__out[15:0];
  assign op_8_53__in1[15:0] = in_107[15:0];
  assign op_8_53__in0[15:0] = in_106[15:0];
  assign op_7_26__in1[15:0] = op_8_53__out[15:0];
  assign op_8_54__in1[15:0] = in_109[15:0];
  assign op_8_54__in0[15:0] = in_108[15:0];
  assign op_7_27__in0[15:0] = op_8_54__out[15:0];
  assign op_8_55__in1[15:0] = in_111[15:0];
  assign op_8_55__in0[15:0] = in_110[15:0];
  assign op_7_27__in1[15:0] = op_8_55__out[15:0];
  assign op_8_56__in1[15:0] = in_113[15:0];
  assign op_8_56__in0[15:0] = in_112[15:0];
  assign op_7_28__in0[15:0] = op_8_56__out[15:0];
  assign op_8_57__in1[15:0] = in_115[15:0];
  assign op_8_57__in0[15:0] = in_114[15:0];
  assign op_7_28__in1[15:0] = op_8_57__out[15:0];
  assign op_8_58__in1[15:0] = in_117[15:0];
  assign op_8_58__in0[15:0] = in_116[15:0];
  assign op_7_29__in0[15:0] = op_8_58__out[15:0];
  assign op_8_59__in1[15:0] = in_119[15:0];
  assign op_8_59__in0[15:0] = in_118[15:0];
  assign op_7_29__in1[15:0] = op_8_59__out[15:0];
  assign op_8_60__in1[15:0] = in_121[15:0];
  assign op_8_60__in0[15:0] = in_120[15:0];
  assign op_7_30__in0[15:0] = op_8_60__out[15:0];
  assign op_8_61__in1[15:0] = in_123[15:0];
  assign op_8_61__in0[15:0] = in_122[15:0];
  assign op_7_30__in1[15:0] = op_8_61__out[15:0];
  assign op_8_62__in1[15:0] = in_125[15:0];
  assign op_8_62__in0[15:0] = in_124[15:0];
  assign op_7_31__in0[15:0] = op_8_62__out[15:0];
  assign op_8_63__in1[15:0] = in_127[15:0];
  assign op_8_63__in0[15:0] = in_126[15:0];
  assign op_7_31__in1[15:0] = op_8_63__out[15:0];
  assign op_8_64__in1[15:0] = in_129[15:0];
  assign op_8_64__in0[15:0] = in_128[15:0];
  assign op_7_32__in0[15:0] = op_8_64__out[15:0];
  assign op_8_65__in1[15:0] = in_131[15:0];
  assign op_8_65__in0[15:0] = in_130[15:0];
  assign op_7_32__in1[15:0] = op_8_65__out[15:0];
  assign op_8_66__in1[15:0] = in_133[15:0];
  assign op_8_66__in0[15:0] = in_132[15:0];
  assign op_7_33__in0[15:0] = op_8_66__out[15:0];
  assign op_8_67__in1[15:0] = in_135[15:0];
  assign op_8_67__in0[15:0] = in_134[15:0];
  assign op_7_33__in1[15:0] = op_8_67__out[15:0];
  assign op_8_68__in1[15:0] = in_137[15:0];
  assign op_8_68__in0[15:0] = in_136[15:0];
  assign op_7_34__in0[15:0] = op_8_68__out[15:0];
  assign op_8_69__in1[15:0] = in_139[15:0];
  assign op_8_69__in0[15:0] = in_138[15:0];
  assign op_7_34__in1[15:0] = op_8_69__out[15:0];
  assign op_8_70__in1[15:0] = in_141[15:0];
  assign op_8_70__in0[15:0] = in_140[15:0];
  assign op_7_35__in0[15:0] = op_8_70__out[15:0];
  assign op_8_71__in1[15:0] = in_143[15:0];
  assign op_8_71__in0[15:0] = in_142[15:0];
  assign op_7_35__in1[15:0] = op_8_71__out[15:0];
  assign op_8_72__in1[15:0] = in_145[15:0];
  assign op_8_72__in0[15:0] = in_144[15:0];
  assign op_7_36__in0[15:0] = op_8_72__out[15:0];
  assign op_8_73__in1[15:0] = in_147[15:0];
  assign op_8_73__in0[15:0] = in_146[15:0];
  assign op_7_36__in1[15:0] = op_8_73__out[15:0];
  assign op_8_74__in1[15:0] = in_149[15:0];
  assign op_8_74__in0[15:0] = in_148[15:0];
  assign op_7_37__in0[15:0] = op_8_74__out[15:0];
  assign op_8_75__in1[15:0] = in_151[15:0];
  assign op_8_75__in0[15:0] = in_150[15:0];
  assign op_7_37__in1[15:0] = op_8_75__out[15:0];
  assign op_8_76__in1[15:0] = in_153[15:0];
  assign op_8_76__in0[15:0] = in_152[15:0];
  assign op_7_38__in0[15:0] = op_8_76__out[15:0];
  assign op_8_77__in1[15:0] = in_155[15:0];
  assign op_8_77__in0[15:0] = in_154[15:0];
  assign op_7_38__in1[15:0] = op_8_77__out[15:0];
  assign op_8_78__in1[15:0] = in_157[15:0];
  assign op_8_78__in0[15:0] = in_156[15:0];
  assign op_7_39__in0[15:0] = op_8_78__out[15:0];
  assign op_8_79__in1[15:0] = in_159[15:0];
  assign op_8_79__in0[15:0] = in_158[15:0];
  assign op_7_39__in1[15:0] = op_8_79__out[15:0];
  assign op_8_80__in1[15:0] = in_161[15:0];
  assign op_8_80__in0[15:0] = in_160[15:0];
  assign op_7_40__in0[15:0] = op_8_80__out[15:0];
  assign op_8_81__in1[15:0] = in_163[15:0];
  assign op_8_81__in0[15:0] = in_162[15:0];
  assign op_7_40__in1[15:0] = op_8_81__out[15:0];
  assign op_8_82__in1[15:0] = in_165[15:0];
  assign op_8_82__in0[15:0] = in_164[15:0];
  assign op_7_41__in0[15:0] = op_8_82__out[15:0];
  assign op_8_83__in1[15:0] = in_167[15:0];
  assign op_8_83__in0[15:0] = in_166[15:0];
  assign op_7_41__in1[15:0] = op_8_83__out[15:0];
  assign op_8_84__in1[15:0] = in_169[15:0];
  assign op_8_84__in0[15:0] = in_168[15:0];
  assign op_7_42__in0[15:0] = op_8_84__out[15:0];
  assign op_8_85__in1[15:0] = in_171[15:0];
  assign op_8_85__in0[15:0] = in_170[15:0];
  assign op_7_42__in1[15:0] = op_8_85__out[15:0];
  assign op_8_86__in1[15:0] = in_173[15:0];
  assign op_8_86__in0[15:0] = in_172[15:0];
  assign op_7_43__in0[15:0] = op_8_86__out[15:0];
  assign op_8_87__in1[15:0] = in_175[15:0];
  assign op_8_87__in0[15:0] = in_174[15:0];
  assign op_7_43__in1[15:0] = op_8_87__out[15:0];
  assign op_8_88__in1[15:0] = in_177[15:0];
  assign op_8_88__in0[15:0] = in_176[15:0];
  assign op_7_44__in0[15:0] = op_8_88__out[15:0];
  assign op_8_89__in1[15:0] = in_179[15:0];
  assign op_8_89__in0[15:0] = in_178[15:0];
  assign op_7_44__in1[15:0] = op_8_89__out[15:0];
  assign op_8_90__in1[15:0] = in_181[15:0];
  assign op_8_90__in0[15:0] = in_180[15:0];
  assign op_7_45__in0[15:0] = op_8_90__out[15:0];
  assign op_8_91__in1[15:0] = in_183[15:0];
  assign op_8_91__in0[15:0] = in_182[15:0];
  assign op_7_45__in1[15:0] = op_8_91__out[15:0];
  assign op_8_92__in1[15:0] = in_185[15:0];
  assign op_8_92__in0[15:0] = in_184[15:0];
  assign op_7_46__in0[15:0] = op_8_92__out[15:0];
  assign op_8_93__in1[15:0] = in_187[15:0];
  assign op_8_93__in0[15:0] = in_186[15:0];
  assign op_7_46__in1[15:0] = op_8_93__out[15:0];
  assign op_8_94__in1[15:0] = in_189[15:0];
  assign op_8_94__in0[15:0] = in_188[15:0];
  assign op_7_47__in0[15:0] = op_8_94__out[15:0];
  assign op_8_95__in1[15:0] = in_191[15:0];
  assign op_8_95__in0[15:0] = in_190[15:0];
  assign op_7_47__in1[15:0] = op_8_95__out[15:0];
  assign op_8_96__in1[15:0] = in_193[15:0];
  assign op_8_96__in0[15:0] = in_192[15:0];
  assign op_7_48__in0[15:0] = op_8_96__out[15:0];
  assign op_8_97__in1[15:0] = in_195[15:0];
  assign op_8_97__in0[15:0] = in_194[15:0];
  assign op_7_48__in1[15:0] = op_8_97__out[15:0];
  assign op_8_98__in1[15:0] = in_197[15:0];
  assign op_8_98__in0[15:0] = in_196[15:0];
  assign op_7_49__in0[15:0] = op_8_98__out[15:0];
  assign op_8_99__in1[15:0] = in_199[15:0];
  assign op_8_99__in0[15:0] = in_198[15:0];
  assign op_7_49__in1[15:0] = op_8_99__out[15:0];
  assign op_8_100__in1[15:0] = in_201[15:0];
  assign op_8_100__in0[15:0] = in_200[15:0];
  assign op_7_50__in0[15:0] = op_8_100__out[15:0];
  assign op_8_101__in1[15:0] = in_203[15:0];
  assign op_8_101__in0[15:0] = in_202[15:0];
  assign op_7_50__in1[15:0] = op_8_101__out[15:0];
  assign op_8_102__in1[15:0] = in_205[15:0];
  assign op_8_102__in0[15:0] = in_204[15:0];
  assign op_7_51__in0[15:0] = op_8_102__out[15:0];
  assign op_8_103__in1[15:0] = in_207[15:0];
  assign op_8_103__in0[15:0] = in_206[15:0];
  assign op_7_51__in1[15:0] = op_8_103__out[15:0];
  assign op_8_104__in1[15:0] = in_209[15:0];
  assign op_8_104__in0[15:0] = in_208[15:0];
  assign op_7_52__in0[15:0] = op_8_104__out[15:0];
  assign op_8_105__in1[15:0] = in_211[15:0];
  assign op_8_105__in0[15:0] = in_210[15:0];
  assign op_7_52__in1[15:0] = op_8_105__out[15:0];
  assign op_8_106__in1[15:0] = in_213[15:0];
  assign op_8_106__in0[15:0] = in_212[15:0];
  assign op_7_53__in0[15:0] = op_8_106__out[15:0];
  assign op_8_107__in1[15:0] = in_215[15:0];
  assign op_8_107__in0[15:0] = in_214[15:0];
  assign op_7_53__in1[15:0] = op_8_107__out[15:0];
  assign op_8_108__in1[15:0] = in_217[15:0];
  assign op_8_108__in0[15:0] = in_216[15:0];
  assign op_7_54__in0[15:0] = op_8_108__out[15:0];
  assign op_8_109__in1[15:0] = in_219[15:0];
  assign op_8_109__in0[15:0] = in_218[15:0];
  assign op_7_54__in1[15:0] = op_8_109__out[15:0];
  assign op_8_110__in1[15:0] = in_221[15:0];
  assign op_8_110__in0[15:0] = in_220[15:0];
  assign op_7_55__in0[15:0] = op_8_110__out[15:0];
  assign op_8_111__in1[15:0] = in_223[15:0];
  assign op_8_111__in0[15:0] = in_222[15:0];
  assign op_7_55__in1[15:0] = op_8_111__out[15:0];
  assign op_8_112__in1[15:0] = in_225[15:0];
  assign op_8_112__in0[15:0] = in_224[15:0];
  assign op_7_56__in0[15:0] = op_8_112__out[15:0];
  assign op_8_113__in1[15:0] = in_227[15:0];
  assign op_8_113__in0[15:0] = in_226[15:0];
  assign op_7_56__in1[15:0] = op_8_113__out[15:0];
  assign op_8_114__in1[15:0] = in_229[15:0];
  assign op_8_114__in0[15:0] = in_228[15:0];
  assign op_7_57__in0[15:0] = op_8_114__out[15:0];
  assign op_8_115__in1[15:0] = in_231[15:0];
  assign op_8_115__in0[15:0] = in_230[15:0];
  assign op_7_57__in1[15:0] = op_8_115__out[15:0];
  assign op_8_116__in1[15:0] = in_233[15:0];
  assign op_8_116__in0[15:0] = in_232[15:0];
  assign op_7_58__in0[15:0] = op_8_116__out[15:0];
  assign op_8_117__in1[15:0] = in_235[15:0];
  assign op_8_117__in0[15:0] = in_234[15:0];
  assign op_7_58__in1[15:0] = op_8_117__out[15:0];
  assign op_8_118__in1[15:0] = in_237[15:0];
  assign op_8_118__in0[15:0] = in_236[15:0];
  assign op_7_59__in0[15:0] = op_8_118__out[15:0];
  assign op_8_119__in1[15:0] = in_239[15:0];
  assign op_8_119__in0[15:0] = in_238[15:0];
  assign op_7_59__in1[15:0] = op_8_119__out[15:0];
  assign op_8_120__in1[15:0] = in_241[15:0];
  assign op_8_120__in0[15:0] = in_240[15:0];
  assign op_7_60__in0[15:0] = op_8_120__out[15:0];
  assign op_8_121__in1[15:0] = in_243[15:0];
  assign op_8_121__in0[15:0] = in_242[15:0];
  assign op_7_60__in1[15:0] = op_8_121__out[15:0];
  assign op_8_122__in1[15:0] = in_245[15:0];
  assign op_8_122__in0[15:0] = in_244[15:0];
  assign op_7_61__in0[15:0] = op_8_122__out[15:0];
  assign op_8_123__in1[15:0] = in_247[15:0];
  assign op_8_123__in0[15:0] = in_246[15:0];
  assign op_7_61__in1[15:0] = op_8_123__out[15:0];
  assign op_8_124__in1[15:0] = in_249[15:0];
  assign op_8_124__in0[15:0] = in_248[15:0];
  assign op_7_62__in0[15:0] = op_8_124__out[15:0];
  assign op_8_125__in1[15:0] = in_251[15:0];
  assign op_8_125__in0[15:0] = in_250[15:0];
  assign op_7_62__in1[15:0] = op_8_125__out[15:0];
  assign op_8_126__in1[15:0] = in_253[15:0];
  assign op_8_126__in0[15:0] = in_252[15:0];
  assign op_7_63__in0[15:0] = op_8_126__out[15:0];
  assign op_8_127__in1[15:0] = in_255[15:0];
  assign op_8_127__in0[15:0] = in_254[15:0];
  assign op_7_63__in1[15:0] = op_8_127__out[15:0];
  assign op_8_128__in1[15:0] = in_257[15:0];
  assign op_8_128__in0[15:0] = in_256[15:0];
  assign op_7_64__in0[15:0] = op_8_128__out[15:0];
  assign op_8_129__in1[15:0] = in_259[15:0];
  assign op_8_129__in0[15:0] = in_258[15:0];
  assign op_7_64__in1[15:0] = op_8_129__out[15:0];
  assign op_8_130__in1[15:0] = in_261[15:0];
  assign op_8_130__in0[15:0] = in_260[15:0];
  assign op_7_65__in0[15:0] = op_8_130__out[15:0];
  assign op_8_131__in1[15:0] = in_263[15:0];
  assign op_8_131__in0[15:0] = in_262[15:0];
  assign op_7_65__in1[15:0] = op_8_131__out[15:0];
  assign op_8_132__in1[15:0] = in_265[15:0];
  assign op_8_132__in0[15:0] = in_264[15:0];
  assign op_7_66__in0[15:0] = op_8_132__out[15:0];
  assign op_8_133__in1[15:0] = in_267[15:0];
  assign op_8_133__in0[15:0] = in_266[15:0];
  assign op_7_66__in1[15:0] = op_8_133__out[15:0];
  assign op_8_134__in1[15:0] = in_269[15:0];
  assign op_8_134__in0[15:0] = in_268[15:0];
  assign op_7_67__in0[15:0] = op_8_134__out[15:0];
  assign op_8_135__in1[15:0] = in_271[15:0];
  assign op_8_135__in0[15:0] = in_270[15:0];
  assign op_7_67__in1[15:0] = op_8_135__out[15:0];
  assign op_8_136__in1[15:0] = in_273[15:0];
  assign op_8_136__in0[15:0] = in_272[15:0];
  assign op_7_68__in0[15:0] = op_8_136__out[15:0];
  assign op_8_137__in1[15:0] = in_275[15:0];
  assign op_8_137__in0[15:0] = in_274[15:0];
  assign op_7_68__in1[15:0] = op_8_137__out[15:0];
  assign op_8_138__in1[15:0] = in_277[15:0];
  assign op_8_138__in0[15:0] = in_276[15:0];
  assign op_7_69__in0[15:0] = op_8_138__out[15:0];
  assign op_8_139__in1[15:0] = in_279[15:0];
  assign op_8_139__in0[15:0] = in_278[15:0];
  assign op_7_69__in1[15:0] = op_8_139__out[15:0];
  assign op_8_140__in1[15:0] = in_281[15:0];
  assign op_8_140__in0[15:0] = in_280[15:0];
  assign op_7_70__in0[15:0] = op_8_140__out[15:0];
  assign op_8_141__in1[15:0] = in_283[15:0];
  assign op_8_141__in0[15:0] = in_282[15:0];
  assign op_7_70__in1[15:0] = op_8_141__out[15:0];
  assign op_8_142__in1[15:0] = in_285[15:0];
  assign op_8_142__in0[15:0] = in_284[15:0];
  assign op_7_71__in0[15:0] = op_8_142__out[15:0];
  assign op_8_143__in1[15:0] = in_287[15:0];
  assign op_8_143__in0[15:0] = in_286[15:0];
  assign op_7_71__in1[15:0] = op_8_143__out[15:0];
  assign op_8_144__in1[15:0] = in_289[15:0];
  assign op_8_144__in0[15:0] = in_288[15:0];
  assign op_7_72__in0[15:0] = op_8_144__out[15:0];
  assign op_8_145__in1[15:0] = in_291[15:0];
  assign op_8_145__in0[15:0] = in_290[15:0];
  assign op_7_72__in1[15:0] = op_8_145__out[15:0];
  assign op_8_146__in1[15:0] = in_293[15:0];
  assign op_8_146__in0[15:0] = in_292[15:0];
  assign op_7_73__in0[15:0] = op_8_146__out[15:0];
  assign op_8_147__in1[15:0] = in_295[15:0];
  assign op_8_147__in0[15:0] = in_294[15:0];
  assign op_7_73__in1[15:0] = op_8_147__out[15:0];
  assign op_8_148__in1[15:0] = in_297[15:0];
  assign op_8_148__in0[15:0] = in_296[15:0];
  assign op_7_74__in0[15:0] = op_8_148__out[15:0];
  assign op_8_149__in1[15:0] = in_299[15:0];
  assign op_8_149__in0[15:0] = in_298[15:0];
  assign op_7_74__in1[15:0] = op_8_149__out[15:0];
  assign op_8_150__in1[15:0] = in_301[15:0];
  assign op_8_150__in0[15:0] = in_300[15:0];
  assign op_7_75__in0[15:0] = op_8_150__out[15:0];
  assign op_8_151__in1[15:0] = in_303[15:0];
  assign op_8_151__in0[15:0] = in_302[15:0];
  assign op_7_75__in1[15:0] = op_8_151__out[15:0];
  assign op_8_152__in1[15:0] = in_305[15:0];
  assign op_8_152__in0[15:0] = in_304[15:0];
  assign op_7_76__in0[15:0] = op_8_152__out[15:0];
  assign op_8_154__in1[15:0] = in_309[15:0];
  assign op_8_154__in0[15:0] = in_308[15:0];
  assign op_7_77__in0[15:0] = op_8_154__out[15:0];
  assign op_8_155__in1[15:0] = in_311[15:0];
  assign op_8_155__in0[15:0] = in_310[15:0];
  assign op_7_77__in1[15:0] = op_8_155__out[15:0];
  assign op_8_156__in1[15:0] = in_313[15:0];
  assign op_8_156__in0[15:0] = in_312[15:0];
  assign op_7_78__in0[15:0] = op_8_156__out[15:0];
  assign op_8_157__in1[15:0] = in_315[15:0];
  assign op_8_157__in0[15:0] = in_314[15:0];
  assign op_7_78__in1[15:0] = op_8_157__out[15:0];
  assign op_8_158__in1[15:0] = in_317[15:0];
  assign op_8_158__in0[15:0] = in_316[15:0];
  assign op_7_79__in0[15:0] = op_8_158__out[15:0];
  assign op_8_159__in1[15:0] = in_319[15:0];
  assign op_8_159__in0[15:0] = in_318[15:0];
  assign op_7_79__in1[15:0] = op_8_159__out[15:0];
  assign op_8_160__in1[15:0] = in_321[15:0];
  assign op_8_160__in0[15:0] = in_320[15:0];
  assign op_7_80__in0[15:0] = op_8_160__out[15:0];
  assign op_8_161__in1[15:0] = in_323[15:0];
  assign op_8_161__in0[15:0] = in_322[15:0];
  assign op_7_80__in1[15:0] = op_8_161__out[15:0];
  assign op_8_162__in1[15:0] = in_325[15:0];
  assign op_8_162__in0[15:0] = in_324[15:0];
  assign op_7_81__in0[15:0] = op_8_162__out[15:0];
  assign op_8_163__in1[15:0] = in_327[15:0];
  assign op_8_163__in0[15:0] = in_326[15:0];
  assign op_7_81__in1[15:0] = op_8_163__out[15:0];
  assign op_8_164__in1[15:0] = in_329[15:0];
  assign op_8_164__in0[15:0] = in_328[15:0];
  assign op_7_82__in0[15:0] = op_8_164__out[15:0];
  assign op_8_165__in1[15:0] = in_331[15:0];
  assign op_8_165__in0[15:0] = in_330[15:0];
  assign op_7_82__in1[15:0] = op_8_165__out[15:0];
  assign op_8_166__in1[15:0] = in_333[15:0];
  assign op_8_166__in0[15:0] = in_332[15:0];
  assign op_7_83__in0[15:0] = op_8_166__out[15:0];
  assign op_8_167__in1[15:0] = in_335[15:0];
  assign op_8_167__in0[15:0] = in_334[15:0];
  assign op_7_83__in1[15:0] = op_8_167__out[15:0];
  assign op_8_168__in1[15:0] = in_337[15:0];
  assign op_8_168__in0[15:0] = in_336[15:0];
  assign op_7_84__in0[15:0] = op_8_168__out[15:0];
  assign op_8_169__in1[15:0] = in_339[15:0];
  assign op_8_169__in0[15:0] = in_338[15:0];
  assign op_7_84__in1[15:0] = op_8_169__out[15:0];
  assign op_8_170__in1[15:0] = in_341[15:0];
  assign op_8_170__in0[15:0] = in_340[15:0];
  assign op_7_85__in0[15:0] = op_8_170__out[15:0];
  assign op_8_171__in1[15:0] = in_343[15:0];
  assign op_8_171__in0[15:0] = in_342[15:0];
  assign op_7_85__in1[15:0] = op_8_171__out[15:0];
  assign op_8_172__in1[15:0] = in_345[15:0];
  assign op_8_172__in0[15:0] = in_344[15:0];
  assign op_7_86__in0[15:0] = op_8_172__out[15:0];
  assign op_8_173__in1[15:0] = in_347[15:0];
  assign op_8_173__in0[15:0] = in_346[15:0];
  assign op_7_86__in1[15:0] = op_8_173__out[15:0];
  assign op_8_174__in1[15:0] = in_349[15:0];
  assign op_8_174__in0[15:0] = in_348[15:0];
  assign op_7_87__in0[15:0] = op_8_174__out[15:0];
  assign op_8_175__in1[15:0] = in_351[15:0];
  assign op_8_175__in0[15:0] = in_350[15:0];
  assign op_7_87__in1[15:0] = op_8_175__out[15:0];
  assign op_8_176__in1[15:0] = in_353[15:0];
  assign op_8_176__in0[15:0] = in_352[15:0];
  assign op_7_88__in0[15:0] = op_8_176__out[15:0];
  assign op_8_177__in1[15:0] = in_355[15:0];
  assign op_8_177__in0[15:0] = in_354[15:0];
  assign op_7_88__in1[15:0] = op_8_177__out[15:0];
  assign op_8_178__in1[15:0] = in_357[15:0];
  assign op_8_178__in0[15:0] = in_356[15:0];
  assign op_7_89__in0[15:0] = op_8_178__out[15:0];
  assign op_8_179__in1[15:0] = in_359[15:0];
  assign op_8_179__in0[15:0] = in_358[15:0];
  assign op_7_89__in1[15:0] = op_8_179__out[15:0];
  assign op_8_180__in1[15:0] = in_361[15:0];
  assign op_8_180__in0[15:0] = in_360[15:0];
  assign op_7_90__in0[15:0] = op_8_180__out[15:0];
  assign op_8_181__in1[15:0] = in_363[15:0];
  assign op_8_181__in0[15:0] = in_362[15:0];
  assign op_7_90__in1[15:0] = op_8_181__out[15:0];
  assign op_8_182__in1[15:0] = in_365[15:0];
  assign op_8_182__in0[15:0] = in_364[15:0];
  assign op_7_91__in0[15:0] = op_8_182__out[15:0];
  assign op_8_183__in1[15:0] = in_367[15:0];
  assign op_8_183__in0[15:0] = in_366[15:0];
  assign op_7_91__in1[15:0] = op_8_183__out[15:0];
  assign op_8_184__in1[15:0] = in_369[15:0];
  assign op_8_184__in0[15:0] = in_368[15:0];
  assign op_7_92__in0[15:0] = op_8_184__out[15:0];
  assign op_8_185__in1[15:0] = in_371[15:0];
  assign op_8_185__in0[15:0] = in_370[15:0];
  assign op_7_92__in1[15:0] = op_8_185__out[15:0];
  assign op_8_186__in1[15:0] = in_373[15:0];
  assign op_8_186__in0[15:0] = in_372[15:0];
  assign op_7_93__in0[15:0] = op_8_186__out[15:0];
  assign op_8_187__in1[15:0] = in_375[15:0];
  assign op_8_187__in0[15:0] = in_374[15:0];
  assign op_7_93__in1[15:0] = op_8_187__out[15:0];
  assign op_8_188__in1[15:0] = in_377[15:0];
  assign op_8_188__in0[15:0] = in_376[15:0];
  assign op_7_94__in0[15:0] = op_8_188__out[15:0];
  assign op_8_189__in1[15:0] = in_379[15:0];
  assign op_8_189__in0[15:0] = in_378[15:0];
  assign op_7_94__in1[15:0] = op_8_189__out[15:0];
  assign op_8_190__in1[15:0] = in_381[15:0];
  assign op_8_190__in0[15:0] = in_380[15:0];
  assign op_7_95__in0[15:0] = op_8_190__out[15:0];
  assign op_8_191__in1[15:0] = in_383[15:0];
  assign op_8_191__in0[15:0] = in_382[15:0];
  assign op_7_95__in1[15:0] = op_8_191__out[15:0];
  assign op_8_192__in1[15:0] = in_385[15:0];
  assign op_8_192__in0[15:0] = in_384[15:0];
  assign op_7_96__in0[15:0] = op_8_192__out[15:0];
  assign op_8_193__in1[15:0] = in_387[15:0];
  assign op_8_193__in0[15:0] = in_386[15:0];
  assign op_7_96__in1[15:0] = op_8_193__out[15:0];
  assign op_8_194__in1[15:0] = in_389[15:0];
  assign op_8_194__in0[15:0] = in_388[15:0];
  assign op_7_97__in0[15:0] = op_8_194__out[15:0];
  assign op_8_195__in1[15:0] = in_391[15:0];
  assign op_8_195__in0[15:0] = in_390[15:0];
  assign op_7_97__in1[15:0] = op_8_195__out[15:0];
  assign op_8_196__in1[15:0] = in_393[15:0];
  assign op_8_196__in0[15:0] = in_392[15:0];
  assign op_7_98__in0[15:0] = op_8_196__out[15:0];
  assign op_8_197__in1[15:0] = in_395[15:0];
  assign op_8_197__in0[15:0] = in_394[15:0];
  assign op_7_98__in1[15:0] = op_8_197__out[15:0];
  assign op_8_198__in1[15:0] = in_397[15:0];
  assign op_8_198__in0[15:0] = in_396[15:0];
  assign op_7_99__in0[15:0] = op_8_198__out[15:0];
  assign op_8_199__in1[15:0] = in_399[15:0];
  assign op_8_199__in0[15:0] = in_398[15:0];
  assign op_7_99__in1[15:0] = op_8_199__out[15:0];
  assign op_8_200__in1[15:0] = in_401[15:0];
  assign op_8_200__in0[15:0] = in_400[15:0];
  assign op_7_100__in0[15:0] = op_8_200__out[15:0];
  assign op_8_201__in1[15:0] = in_403[15:0];
  assign op_8_201__in0[15:0] = in_402[15:0];
  assign op_7_100__in1[15:0] = op_8_201__out[15:0];
  assign op_8_202__in1[15:0] = in_405[15:0];
  assign op_8_202__in0[15:0] = in_404[15:0];
  assign op_7_101__in0[15:0] = op_8_202__out[15:0];
  assign op_8_203__in1[15:0] = in_407[15:0];
  assign op_8_203__in0[15:0] = in_406[15:0];
  assign op_7_101__in1[15:0] = op_8_203__out[15:0];
  assign op_8_204__in1[15:0] = in_409[15:0];
  assign op_8_204__in0[15:0] = in_408[15:0];
  assign op_7_102__in0[15:0] = op_8_204__out[15:0];
  assign op_8_205__in1[15:0] = in_411[15:0];
  assign op_8_205__in0[15:0] = in_410[15:0];
  assign op_7_102__in1[15:0] = op_8_205__out[15:0];
  assign op_8_206__in1[15:0] = in_413[15:0];
  assign op_8_206__in0[15:0] = in_412[15:0];
  assign op_7_103__in0[15:0] = op_8_206__out[15:0];
  assign op_8_207__in1[15:0] = in_415[15:0];
  assign op_8_207__in0[15:0] = in_414[15:0];
  assign op_7_103__in1[15:0] = op_8_207__out[15:0];
  assign op_8_208__in1[15:0] = in_417[15:0];
  assign op_8_208__in0[15:0] = in_416[15:0];
  assign op_7_104__in0[15:0] = op_8_208__out[15:0];
  assign op_8_209__in1[15:0] = in_419[15:0];
  assign op_8_209__in0[15:0] = in_418[15:0];
  assign op_7_104__in1[15:0] = op_8_209__out[15:0];
  assign op_8_210__in1[15:0] = in_421[15:0];
  assign op_8_210__in0[15:0] = in_420[15:0];
  assign op_7_105__in0[15:0] = op_8_210__out[15:0];
  assign op_8_211__in1[15:0] = in_423[15:0];
  assign op_8_211__in0[15:0] = in_422[15:0];
  assign op_7_105__in1[15:0] = op_8_211__out[15:0];
  assign op_8_212__in1[15:0] = in_425[15:0];
  assign op_8_212__in0[15:0] = in_424[15:0];
  assign op_7_106__in0[15:0] = op_8_212__out[15:0];
  assign op_8_213__in1[15:0] = in_427[15:0];
  assign op_8_213__in0[15:0] = in_426[15:0];
  assign op_7_106__in1[15:0] = op_8_213__out[15:0];
  assign op_8_214__in1[15:0] = in_429[15:0];
  assign op_8_214__in0[15:0] = in_428[15:0];
  assign op_7_107__in0[15:0] = op_8_214__out[15:0];
  assign op_8_215__in1[15:0] = in_431[15:0];
  assign op_8_215__in0[15:0] = in_430[15:0];
  assign op_7_107__in1[15:0] = op_8_215__out[15:0];
  assign op_8_216__in1[15:0] = in_433[15:0];
  assign op_8_216__in0[15:0] = in_432[15:0];
  assign op_7_108__in0[15:0] = op_8_216__out[15:0];
  assign op_8_217__in1[15:0] = in_435[15:0];
  assign op_8_217__in0[15:0] = in_434[15:0];
  assign op_7_108__in1[15:0] = op_8_217__out[15:0];
  assign op_8_218__in1[15:0] = in_437[15:0];
  assign op_8_218__in0[15:0] = in_436[15:0];
  assign op_7_109__in0[15:0] = op_8_218__out[15:0];
  assign op_8_219__in1[15:0] = in_439[15:0];
  assign op_8_219__in0[15:0] = in_438[15:0];
  assign op_7_109__in1[15:0] = op_8_219__out[15:0];
  assign op_8_220__in1[15:0] = in_441[15:0];
  assign op_8_220__in0[15:0] = in_440[15:0];
  assign op_7_110__in0[15:0] = op_8_220__out[15:0];
  assign op_8_221__in1[15:0] = in_443[15:0];
  assign op_8_221__in0[15:0] = in_442[15:0];
  assign op_7_110__in1[15:0] = op_8_221__out[15:0];
  assign op_8_222__in1[15:0] = in_445[15:0];
  assign op_8_222__in0[15:0] = in_444[15:0];
  assign op_7_111__in0[15:0] = op_8_222__out[15:0];
  assign op_8_223__in1[15:0] = in_447[15:0];
  assign op_8_223__in0[15:0] = in_446[15:0];
  assign op_7_111__in1[15:0] = op_8_223__out[15:0];
  assign op_8_224__in1[15:0] = in_449[15:0];
  assign op_8_224__in0[15:0] = in_448[15:0];
  assign op_7_112__in0[15:0] = op_8_224__out[15:0];
  assign op_8_225__in1[15:0] = in_451[15:0];
  assign op_8_225__in0[15:0] = in_450[15:0];
  assign op_7_112__in1[15:0] = op_8_225__out[15:0];
  assign op_8_226__in1[15:0] = in_453[15:0];
  assign op_8_226__in0[15:0] = in_452[15:0];
  assign op_7_113__in0[15:0] = op_8_226__out[15:0];
  assign op_8_227__in1[15:0] = in_455[15:0];
  assign op_8_227__in0[15:0] = in_454[15:0];
  assign op_7_113__in1[15:0] = op_8_227__out[15:0];
  assign op_8_228__in1[15:0] = in_457[15:0];
  assign op_8_228__in0[15:0] = in_456[15:0];
  assign op_7_114__in0[15:0] = op_8_228__out[15:0];
  assign op_8_229__in1[15:0] = in_459[15:0];
  assign op_8_229__in0[15:0] = in_458[15:0];
  assign op_7_114__in1[15:0] = op_8_229__out[15:0];
  assign op_8_230__in1[15:0] = in_461[15:0];
  assign op_8_230__in0[15:0] = in_460[15:0];
  assign op_7_115__in0[15:0] = op_8_230__out[15:0];
  assign op_8_231__in1[15:0] = in_463[15:0];
  assign op_8_231__in0[15:0] = in_462[15:0];
  assign op_7_115__in1[15:0] = op_8_231__out[15:0];
  assign op_8_232__in1[15:0] = in_465[15:0];
  assign op_8_232__in0[15:0] = in_464[15:0];
  assign op_7_116__in0[15:0] = op_8_232__out[15:0];
  assign op_8_233__in1[15:0] = in_467[15:0];
  assign op_8_233__in0[15:0] = in_466[15:0];
  assign op_7_116__in1[15:0] = op_8_233__out[15:0];
  assign op_8_234__in1[15:0] = in_469[15:0];
  assign op_8_234__in0[15:0] = in_468[15:0];
  assign op_7_117__in0[15:0] = op_8_234__out[15:0];
  assign op_8_235__in1[15:0] = in_471[15:0];
  assign op_8_235__in0[15:0] = in_470[15:0];
  assign op_7_117__in1[15:0] = op_8_235__out[15:0];
  assign op_8_236__in1[15:0] = in_473[15:0];
  assign op_8_236__in0[15:0] = in_472[15:0];
  assign op_7_118__in0[15:0] = op_8_236__out[15:0];
  assign op_8_237__in1[15:0] = in_475[15:0];
  assign op_8_237__in0[15:0] = in_474[15:0];
  assign op_7_118__in1[15:0] = op_8_237__out[15:0];
  assign op_8_238__in1[15:0] = in_477[15:0];
  assign op_8_238__in0[15:0] = in_476[15:0];
  assign op_7_119__in0[15:0] = op_8_238__out[15:0];
  assign op_8_239__in1[15:0] = in_479[15:0];
  assign op_8_239__in0[15:0] = in_478[15:0];
  assign op_7_119__in1[15:0] = op_8_239__out[15:0];
  assign op_8_240__in1[15:0] = in_481[15:0];
  assign op_8_240__in0[15:0] = in_480[15:0];
  assign op_7_120__in0[15:0] = op_8_240__out[15:0];
  assign op_8_241__in1[15:0] = in_483[15:0];
  assign op_8_241__in0[15:0] = in_482[15:0];
  assign op_7_120__in1[15:0] = op_8_241__out[15:0];
  assign op_8_242__in1[15:0] = in_485[15:0];
  assign op_8_242__in0[15:0] = in_484[15:0];
  assign op_7_121__in0[15:0] = op_8_242__out[15:0];
  assign op_8_243__in1[15:0] = in_487[15:0];
  assign op_8_243__in0[15:0] = in_486[15:0];
  assign op_7_121__in1[15:0] = op_8_243__out[15:0];
  assign op_8_244__in1[15:0] = in_489[15:0];
  assign op_8_244__in0[15:0] = in_488[15:0];
  assign op_7_122__in0[15:0] = op_8_244__out[15:0];
  assign op_8_245__in1[15:0] = in_491[15:0];
  assign op_8_245__in0[15:0] = in_490[15:0];
  assign op_7_122__in1[15:0] = op_8_245__out[15:0];
  assign op_8_246__in1[15:0] = in_493[15:0];
  assign op_8_246__in0[15:0] = in_492[15:0];
  assign op_7_123__in0[15:0] = op_8_246__out[15:0];
  assign op_8_247__in1[15:0] = in_495[15:0];
  assign op_8_247__in0[15:0] = in_494[15:0];
  assign op_7_123__in1[15:0] = op_8_247__out[15:0];
  assign op_8_248__in1[15:0] = in_497[15:0];
  assign op_8_248__in0[15:0] = in_496[15:0];
  assign op_7_124__in0[15:0] = op_8_248__out[15:0];
  assign op_8_249__in1[15:0] = in_499[15:0];
  assign op_8_249__in0[15:0] = in_498[15:0];
  assign op_7_124__in1[15:0] = op_8_249__out[15:0];
  assign op_8_250__in1[15:0] = in_501[15:0];
  assign op_8_250__in0[15:0] = in_500[15:0];
  assign op_7_125__in0[15:0] = op_8_250__out[15:0];
  assign op_8_251__in1[15:0] = in_503[15:0];
  assign op_8_251__in0[15:0] = in_502[15:0];
  assign op_7_125__in1[15:0] = op_8_251__out[15:0];
  assign op_8_252__in1[15:0] = in_505[15:0];
  assign op_8_252__in0[15:0] = in_504[15:0];
  assign op_7_126__in0[15:0] = op_8_252__out[15:0];
  assign op_8_253__in1[15:0] = in_507[15:0];
  assign op_8_253__in0[15:0] = in_506[15:0];
  assign op_7_126__in1[15:0] = op_8_253__out[15:0];
  assign op_8_254__in1[15:0] = in_509[15:0];
  assign op_8_254__in0[15:0] = in_508[15:0];
  assign op_7_127__in0[15:0] = op_8_254__out[15:0];
  assign op_8_255__in1[15:0] = in_511[15:0];
  assign op_8_255__in0[15:0] = in_510[15:0];
  assign op_7_127__in1[15:0] = op_8_255__out[15:0];

endmodule //reduceParallelPower2Inputs_U2

module reduceParallel_U1 (
  input [15:0] in_data_0,
  input [15:0] in_data_1,
  input [15:0] in_data_10,
  input [15:0] in_data_100,
  input [15:0] in_data_101,
  input [15:0] in_data_102,
  input [15:0] in_data_103,
  input [15:0] in_data_104,
  input [15:0] in_data_105,
  input [15:0] in_data_106,
  input [15:0] in_data_107,
  input [15:0] in_data_108,
  input [15:0] in_data_109,
  input [15:0] in_data_11,
  input [15:0] in_data_110,
  input [15:0] in_data_111,
  input [15:0] in_data_112,
  input [15:0] in_data_113,
  input [15:0] in_data_114,
  input [15:0] in_data_115,
  input [15:0] in_data_116,
  input [15:0] in_data_117,
  input [15:0] in_data_118,
  input [15:0] in_data_119,
  input [15:0] in_data_12,
  input [15:0] in_data_120,
  input [15:0] in_data_121,
  input [15:0] in_data_122,
  input [15:0] in_data_123,
  input [15:0] in_data_124,
  input [15:0] in_data_125,
  input [15:0] in_data_126,
  input [15:0] in_data_127,
  input [15:0] in_data_128,
  input [15:0] in_data_129,
  input [15:0] in_data_13,
  input [15:0] in_data_130,
  input [15:0] in_data_131,
  input [15:0] in_data_132,
  input [15:0] in_data_133,
  input [15:0] in_data_134,
  input [15:0] in_data_135,
  input [15:0] in_data_136,
  input [15:0] in_data_137,
  input [15:0] in_data_138,
  input [15:0] in_data_139,
  input [15:0] in_data_14,
  input [15:0] in_data_140,
  input [15:0] in_data_141,
  input [15:0] in_data_142,
  input [15:0] in_data_143,
  input [15:0] in_data_144,
  input [15:0] in_data_145,
  input [15:0] in_data_146,
  input [15:0] in_data_147,
  input [15:0] in_data_148,
  input [15:0] in_data_149,
  input [15:0] in_data_15,
  input [15:0] in_data_150,
  input [15:0] in_data_151,
  input [15:0] in_data_152,
  input [15:0] in_data_153,
  input [15:0] in_data_154,
  input [15:0] in_data_155,
  input [15:0] in_data_156,
  input [15:0] in_data_157,
  input [15:0] in_data_158,
  input [15:0] in_data_159,
  input [15:0] in_data_16,
  input [15:0] in_data_160,
  input [15:0] in_data_161,
  input [15:0] in_data_162,
  input [15:0] in_data_163,
  input [15:0] in_data_164,
  input [15:0] in_data_165,
  input [15:0] in_data_166,
  input [15:0] in_data_167,
  input [15:0] in_data_168,
  input [15:0] in_data_169,
  input [15:0] in_data_17,
  input [15:0] in_data_170,
  input [15:0] in_data_171,
  input [15:0] in_data_172,
  input [15:0] in_data_173,
  input [15:0] in_data_174,
  input [15:0] in_data_175,
  input [15:0] in_data_176,
  input [15:0] in_data_177,
  input [15:0] in_data_178,
  input [15:0] in_data_179,
  input [15:0] in_data_18,
  input [15:0] in_data_180,
  input [15:0] in_data_181,
  input [15:0] in_data_182,
  input [15:0] in_data_183,
  input [15:0] in_data_184,
  input [15:0] in_data_185,
  input [15:0] in_data_186,
  input [15:0] in_data_187,
  input [15:0] in_data_188,
  input [15:0] in_data_189,
  input [15:0] in_data_19,
  input [15:0] in_data_190,
  input [15:0] in_data_191,
  input [15:0] in_data_192,
  input [15:0] in_data_193,
  input [15:0] in_data_194,
  input [15:0] in_data_195,
  input [15:0] in_data_196,
  input [15:0] in_data_197,
  input [15:0] in_data_198,
  input [15:0] in_data_199,
  input [15:0] in_data_2,
  input [15:0] in_data_20,
  input [15:0] in_data_200,
  input [15:0] in_data_201,
  input [15:0] in_data_202,
  input [15:0] in_data_203,
  input [15:0] in_data_204,
  input [15:0] in_data_205,
  input [15:0] in_data_206,
  input [15:0] in_data_207,
  input [15:0] in_data_208,
  input [15:0] in_data_209,
  input [15:0] in_data_21,
  input [15:0] in_data_210,
  input [15:0] in_data_211,
  input [15:0] in_data_212,
  input [15:0] in_data_213,
  input [15:0] in_data_214,
  input [15:0] in_data_215,
  input [15:0] in_data_216,
  input [15:0] in_data_217,
  input [15:0] in_data_218,
  input [15:0] in_data_219,
  input [15:0] in_data_22,
  input [15:0] in_data_220,
  input [15:0] in_data_221,
  input [15:0] in_data_222,
  input [15:0] in_data_223,
  input [15:0] in_data_224,
  input [15:0] in_data_225,
  input [15:0] in_data_226,
  input [15:0] in_data_227,
  input [15:0] in_data_228,
  input [15:0] in_data_229,
  input [15:0] in_data_23,
  input [15:0] in_data_230,
  input [15:0] in_data_231,
  input [15:0] in_data_232,
  input [15:0] in_data_233,
  input [15:0] in_data_234,
  input [15:0] in_data_235,
  input [15:0] in_data_236,
  input [15:0] in_data_237,
  input [15:0] in_data_238,
  input [15:0] in_data_239,
  input [15:0] in_data_24,
  input [15:0] in_data_240,
  input [15:0] in_data_241,
  input [15:0] in_data_242,
  input [15:0] in_data_243,
  input [15:0] in_data_244,
  input [15:0] in_data_245,
  input [15:0] in_data_246,
  input [15:0] in_data_247,
  input [15:0] in_data_248,
  input [15:0] in_data_249,
  input [15:0] in_data_25,
  input [15:0] in_data_250,
  input [15:0] in_data_251,
  input [15:0] in_data_252,
  input [15:0] in_data_253,
  input [15:0] in_data_254,
  input [15:0] in_data_255,
  input [15:0] in_data_256,
  input [15:0] in_data_257,
  input [15:0] in_data_258,
  input [15:0] in_data_259,
  input [15:0] in_data_26,
  input [15:0] in_data_260,
  input [15:0] in_data_261,
  input [15:0] in_data_262,
  input [15:0] in_data_263,
  input [15:0] in_data_264,
  input [15:0] in_data_265,
  input [15:0] in_data_266,
  input [15:0] in_data_267,
  input [15:0] in_data_268,
  input [15:0] in_data_269,
  input [15:0] in_data_27,
  input [15:0] in_data_270,
  input [15:0] in_data_271,
  input [15:0] in_data_272,
  input [15:0] in_data_273,
  input [15:0] in_data_274,
  input [15:0] in_data_275,
  input [15:0] in_data_276,
  input [15:0] in_data_277,
  input [15:0] in_data_278,
  input [15:0] in_data_279,
  input [15:0] in_data_28,
  input [15:0] in_data_280,
  input [15:0] in_data_281,
  input [15:0] in_data_282,
  input [15:0] in_data_283,
  input [15:0] in_data_284,
  input [15:0] in_data_285,
  input [15:0] in_data_286,
  input [15:0] in_data_287,
  input [15:0] in_data_288,
  input [15:0] in_data_289,
  input [15:0] in_data_29,
  input [15:0] in_data_290,
  input [15:0] in_data_291,
  input [15:0] in_data_292,
  input [15:0] in_data_293,
  input [15:0] in_data_294,
  input [15:0] in_data_295,
  input [15:0] in_data_296,
  input [15:0] in_data_297,
  input [15:0] in_data_298,
  input [15:0] in_data_299,
  input [15:0] in_data_3,
  input [15:0] in_data_30,
  input [15:0] in_data_31,
  input [15:0] in_data_32,
  input [15:0] in_data_33,
  input [15:0] in_data_34,
  input [15:0] in_data_35,
  input [15:0] in_data_36,
  input [15:0] in_data_37,
  input [15:0] in_data_38,
  input [15:0] in_data_39,
  input [15:0] in_data_4,
  input [15:0] in_data_40,
  input [15:0] in_data_41,
  input [15:0] in_data_42,
  input [15:0] in_data_43,
  input [15:0] in_data_44,
  input [15:0] in_data_45,
  input [15:0] in_data_46,
  input [15:0] in_data_47,
  input [15:0] in_data_48,
  input [15:0] in_data_49,
  input [15:0] in_data_5,
  input [15:0] in_data_50,
  input [15:0] in_data_51,
  input [15:0] in_data_52,
  input [15:0] in_data_53,
  input [15:0] in_data_54,
  input [15:0] in_data_55,
  input [15:0] in_data_56,
  input [15:0] in_data_57,
  input [15:0] in_data_58,
  input [15:0] in_data_59,
  input [15:0] in_data_6,
  input [15:0] in_data_60,
  input [15:0] in_data_61,
  input [15:0] in_data_62,
  input [15:0] in_data_63,
  input [15:0] in_data_64,
  input [15:0] in_data_65,
  input [15:0] in_data_66,
  input [15:0] in_data_67,
  input [15:0] in_data_68,
  input [15:0] in_data_69,
  input [15:0] in_data_7,
  input [15:0] in_data_70,
  input [15:0] in_data_71,
  input [15:0] in_data_72,
  input [15:0] in_data_73,
  input [15:0] in_data_74,
  input [15:0] in_data_75,
  input [15:0] in_data_76,
  input [15:0] in_data_77,
  input [15:0] in_data_78,
  input [15:0] in_data_79,
  input [15:0] in_data_8,
  input [15:0] in_data_80,
  input [15:0] in_data_81,
  input [15:0] in_data_82,
  input [15:0] in_data_83,
  input [15:0] in_data_84,
  input [15:0] in_data_85,
  input [15:0] in_data_86,
  input [15:0] in_data_87,
  input [15:0] in_data_88,
  input [15:0] in_data_89,
  input [15:0] in_data_9,
  input [15:0] in_data_90,
  input [15:0] in_data_91,
  input [15:0] in_data_92,
  input [15:0] in_data_93,
  input [15:0] in_data_94,
  input [15:0] in_data_95,
  input [15:0] in_data_96,
  input [15:0] in_data_97,
  input [15:0] in_data_98,
  input [15:0] in_data_99,
  input [15:0] in_identity,
  output [15:0] out
);
  //Wire declarations for instance 'reducer' (Module reduceParallelPower2Inputs_U2)
  wire [15:0] reducer__in_0;
  wire [15:0] reducer__in_1;
  wire [15:0] reducer__in_10;
  wire [15:0] reducer__in_100;
  wire [15:0] reducer__in_101;
  wire [15:0] reducer__in_102;
  wire [15:0] reducer__in_103;
  wire [15:0] reducer__in_104;
  wire [15:0] reducer__in_105;
  wire [15:0] reducer__in_106;
  wire [15:0] reducer__in_107;
  wire [15:0] reducer__in_108;
  wire [15:0] reducer__in_109;
  wire [15:0] reducer__in_11;
  wire [15:0] reducer__in_110;
  wire [15:0] reducer__in_111;
  wire [15:0] reducer__in_112;
  wire [15:0] reducer__in_113;
  wire [15:0] reducer__in_114;
  wire [15:0] reducer__in_115;
  wire [15:0] reducer__in_116;
  wire [15:0] reducer__in_117;
  wire [15:0] reducer__in_118;
  wire [15:0] reducer__in_119;
  wire [15:0] reducer__in_12;
  wire [15:0] reducer__in_120;
  wire [15:0] reducer__in_121;
  wire [15:0] reducer__in_122;
  wire [15:0] reducer__in_123;
  wire [15:0] reducer__in_124;
  wire [15:0] reducer__in_125;
  wire [15:0] reducer__in_126;
  wire [15:0] reducer__in_127;
  wire [15:0] reducer__in_128;
  wire [15:0] reducer__in_129;
  wire [15:0] reducer__in_13;
  wire [15:0] reducer__in_130;
  wire [15:0] reducer__in_131;
  wire [15:0] reducer__in_132;
  wire [15:0] reducer__in_133;
  wire [15:0] reducer__in_134;
  wire [15:0] reducer__in_135;
  wire [15:0] reducer__in_136;
  wire [15:0] reducer__in_137;
  wire [15:0] reducer__in_138;
  wire [15:0] reducer__in_139;
  wire [15:0] reducer__in_14;
  wire [15:0] reducer__in_140;
  wire [15:0] reducer__in_141;
  wire [15:0] reducer__in_142;
  wire [15:0] reducer__in_143;
  wire [15:0] reducer__in_144;
  wire [15:0] reducer__in_145;
  wire [15:0] reducer__in_146;
  wire [15:0] reducer__in_147;
  wire [15:0] reducer__in_148;
  wire [15:0] reducer__in_149;
  wire [15:0] reducer__in_15;
  wire [15:0] reducer__in_150;
  wire [15:0] reducer__in_151;
  wire [15:0] reducer__in_152;
  wire [15:0] reducer__in_153;
  wire [15:0] reducer__in_154;
  wire [15:0] reducer__in_155;
  wire [15:0] reducer__in_156;
  wire [15:0] reducer__in_157;
  wire [15:0] reducer__in_158;
  wire [15:0] reducer__in_159;
  wire [15:0] reducer__in_16;
  wire [15:0] reducer__in_160;
  wire [15:0] reducer__in_161;
  wire [15:0] reducer__in_162;
  wire [15:0] reducer__in_163;
  wire [15:0] reducer__in_164;
  wire [15:0] reducer__in_165;
  wire [15:0] reducer__in_166;
  wire [15:0] reducer__in_167;
  wire [15:0] reducer__in_168;
  wire [15:0] reducer__in_169;
  wire [15:0] reducer__in_17;
  wire [15:0] reducer__in_170;
  wire [15:0] reducer__in_171;
  wire [15:0] reducer__in_172;
  wire [15:0] reducer__in_173;
  wire [15:0] reducer__in_174;
  wire [15:0] reducer__in_175;
  wire [15:0] reducer__in_176;
  wire [15:0] reducer__in_177;
  wire [15:0] reducer__in_178;
  wire [15:0] reducer__in_179;
  wire [15:0] reducer__in_18;
  wire [15:0] reducer__in_180;
  wire [15:0] reducer__in_181;
  wire [15:0] reducer__in_182;
  wire [15:0] reducer__in_183;
  wire [15:0] reducer__in_184;
  wire [15:0] reducer__in_185;
  wire [15:0] reducer__in_186;
  wire [15:0] reducer__in_187;
  wire [15:0] reducer__in_188;
  wire [15:0] reducer__in_189;
  wire [15:0] reducer__in_19;
  wire [15:0] reducer__in_190;
  wire [15:0] reducer__in_191;
  wire [15:0] reducer__in_192;
  wire [15:0] reducer__in_193;
  wire [15:0] reducer__in_194;
  wire [15:0] reducer__in_195;
  wire [15:0] reducer__in_196;
  wire [15:0] reducer__in_197;
  wire [15:0] reducer__in_198;
  wire [15:0] reducer__in_199;
  wire [15:0] reducer__in_2;
  wire [15:0] reducer__in_20;
  wire [15:0] reducer__in_200;
  wire [15:0] reducer__in_201;
  wire [15:0] reducer__in_202;
  wire [15:0] reducer__in_203;
  wire [15:0] reducer__in_204;
  wire [15:0] reducer__in_205;
  wire [15:0] reducer__in_206;
  wire [15:0] reducer__in_207;
  wire [15:0] reducer__in_208;
  wire [15:0] reducer__in_209;
  wire [15:0] reducer__in_21;
  wire [15:0] reducer__in_210;
  wire [15:0] reducer__in_211;
  wire [15:0] reducer__in_212;
  wire [15:0] reducer__in_213;
  wire [15:0] reducer__in_214;
  wire [15:0] reducer__in_215;
  wire [15:0] reducer__in_216;
  wire [15:0] reducer__in_217;
  wire [15:0] reducer__in_218;
  wire [15:0] reducer__in_219;
  wire [15:0] reducer__in_22;
  wire [15:0] reducer__in_220;
  wire [15:0] reducer__in_221;
  wire [15:0] reducer__in_222;
  wire [15:0] reducer__in_223;
  wire [15:0] reducer__in_224;
  wire [15:0] reducer__in_225;
  wire [15:0] reducer__in_226;
  wire [15:0] reducer__in_227;
  wire [15:0] reducer__in_228;
  wire [15:0] reducer__in_229;
  wire [15:0] reducer__in_23;
  wire [15:0] reducer__in_230;
  wire [15:0] reducer__in_231;
  wire [15:0] reducer__in_232;
  wire [15:0] reducer__in_233;
  wire [15:0] reducer__in_234;
  wire [15:0] reducer__in_235;
  wire [15:0] reducer__in_236;
  wire [15:0] reducer__in_237;
  wire [15:0] reducer__in_238;
  wire [15:0] reducer__in_239;
  wire [15:0] reducer__in_24;
  wire [15:0] reducer__in_240;
  wire [15:0] reducer__in_241;
  wire [15:0] reducer__in_242;
  wire [15:0] reducer__in_243;
  wire [15:0] reducer__in_244;
  wire [15:0] reducer__in_245;
  wire [15:0] reducer__in_246;
  wire [15:0] reducer__in_247;
  wire [15:0] reducer__in_248;
  wire [15:0] reducer__in_249;
  wire [15:0] reducer__in_25;
  wire [15:0] reducer__in_250;
  wire [15:0] reducer__in_251;
  wire [15:0] reducer__in_252;
  wire [15:0] reducer__in_253;
  wire [15:0] reducer__in_254;
  wire [15:0] reducer__in_255;
  wire [15:0] reducer__in_256;
  wire [15:0] reducer__in_257;
  wire [15:0] reducer__in_258;
  wire [15:0] reducer__in_259;
  wire [15:0] reducer__in_26;
  wire [15:0] reducer__in_260;
  wire [15:0] reducer__in_261;
  wire [15:0] reducer__in_262;
  wire [15:0] reducer__in_263;
  wire [15:0] reducer__in_264;
  wire [15:0] reducer__in_265;
  wire [15:0] reducer__in_266;
  wire [15:0] reducer__in_267;
  wire [15:0] reducer__in_268;
  wire [15:0] reducer__in_269;
  wire [15:0] reducer__in_27;
  wire [15:0] reducer__in_270;
  wire [15:0] reducer__in_271;
  wire [15:0] reducer__in_272;
  wire [15:0] reducer__in_273;
  wire [15:0] reducer__in_274;
  wire [15:0] reducer__in_275;
  wire [15:0] reducer__in_276;
  wire [15:0] reducer__in_277;
  wire [15:0] reducer__in_278;
  wire [15:0] reducer__in_279;
  wire [15:0] reducer__in_28;
  wire [15:0] reducer__in_280;
  wire [15:0] reducer__in_281;
  wire [15:0] reducer__in_282;
  wire [15:0] reducer__in_283;
  wire [15:0] reducer__in_284;
  wire [15:0] reducer__in_285;
  wire [15:0] reducer__in_286;
  wire [15:0] reducer__in_287;
  wire [15:0] reducer__in_288;
  wire [15:0] reducer__in_289;
  wire [15:0] reducer__in_29;
  wire [15:0] reducer__in_290;
  wire [15:0] reducer__in_291;
  wire [15:0] reducer__in_292;
  wire [15:0] reducer__in_293;
  wire [15:0] reducer__in_294;
  wire [15:0] reducer__in_295;
  wire [15:0] reducer__in_296;
  wire [15:0] reducer__in_297;
  wire [15:0] reducer__in_298;
  wire [15:0] reducer__in_299;
  wire [15:0] reducer__in_3;
  wire [15:0] reducer__in_30;
  wire [15:0] reducer__in_300;
  wire [15:0] reducer__in_301;
  wire [15:0] reducer__in_302;
  wire [15:0] reducer__in_303;
  wire [15:0] reducer__in_304;
  wire [15:0] reducer__in_305;
  wire [15:0] reducer__in_306;
  wire [15:0] reducer__in_307;
  wire [15:0] reducer__in_308;
  wire [15:0] reducer__in_309;
  wire [15:0] reducer__in_31;
  wire [15:0] reducer__in_310;
  wire [15:0] reducer__in_311;
  wire [15:0] reducer__in_312;
  wire [15:0] reducer__in_313;
  wire [15:0] reducer__in_314;
  wire [15:0] reducer__in_315;
  wire [15:0] reducer__in_316;
  wire [15:0] reducer__in_317;
  wire [15:0] reducer__in_318;
  wire [15:0] reducer__in_319;
  wire [15:0] reducer__in_32;
  wire [15:0] reducer__in_320;
  wire [15:0] reducer__in_321;
  wire [15:0] reducer__in_322;
  wire [15:0] reducer__in_323;
  wire [15:0] reducer__in_324;
  wire [15:0] reducer__in_325;
  wire [15:0] reducer__in_326;
  wire [15:0] reducer__in_327;
  wire [15:0] reducer__in_328;
  wire [15:0] reducer__in_329;
  wire [15:0] reducer__in_33;
  wire [15:0] reducer__in_330;
  wire [15:0] reducer__in_331;
  wire [15:0] reducer__in_332;
  wire [15:0] reducer__in_333;
  wire [15:0] reducer__in_334;
  wire [15:0] reducer__in_335;
  wire [15:0] reducer__in_336;
  wire [15:0] reducer__in_337;
  wire [15:0] reducer__in_338;
  wire [15:0] reducer__in_339;
  wire [15:0] reducer__in_34;
  wire [15:0] reducer__in_340;
  wire [15:0] reducer__in_341;
  wire [15:0] reducer__in_342;
  wire [15:0] reducer__in_343;
  wire [15:0] reducer__in_344;
  wire [15:0] reducer__in_345;
  wire [15:0] reducer__in_346;
  wire [15:0] reducer__in_347;
  wire [15:0] reducer__in_348;
  wire [15:0] reducer__in_349;
  wire [15:0] reducer__in_35;
  wire [15:0] reducer__in_350;
  wire [15:0] reducer__in_351;
  wire [15:0] reducer__in_352;
  wire [15:0] reducer__in_353;
  wire [15:0] reducer__in_354;
  wire [15:0] reducer__in_355;
  wire [15:0] reducer__in_356;
  wire [15:0] reducer__in_357;
  wire [15:0] reducer__in_358;
  wire [15:0] reducer__in_359;
  wire [15:0] reducer__in_36;
  wire [15:0] reducer__in_360;
  wire [15:0] reducer__in_361;
  wire [15:0] reducer__in_362;
  wire [15:0] reducer__in_363;
  wire [15:0] reducer__in_364;
  wire [15:0] reducer__in_365;
  wire [15:0] reducer__in_366;
  wire [15:0] reducer__in_367;
  wire [15:0] reducer__in_368;
  wire [15:0] reducer__in_369;
  wire [15:0] reducer__in_37;
  wire [15:0] reducer__in_370;
  wire [15:0] reducer__in_371;
  wire [15:0] reducer__in_372;
  wire [15:0] reducer__in_373;
  wire [15:0] reducer__in_374;
  wire [15:0] reducer__in_375;
  wire [15:0] reducer__in_376;
  wire [15:0] reducer__in_377;
  wire [15:0] reducer__in_378;
  wire [15:0] reducer__in_379;
  wire [15:0] reducer__in_38;
  wire [15:0] reducer__in_380;
  wire [15:0] reducer__in_381;
  wire [15:0] reducer__in_382;
  wire [15:0] reducer__in_383;
  wire [15:0] reducer__in_384;
  wire [15:0] reducer__in_385;
  wire [15:0] reducer__in_386;
  wire [15:0] reducer__in_387;
  wire [15:0] reducer__in_388;
  wire [15:0] reducer__in_389;
  wire [15:0] reducer__in_39;
  wire [15:0] reducer__in_390;
  wire [15:0] reducer__in_391;
  wire [15:0] reducer__in_392;
  wire [15:0] reducer__in_393;
  wire [15:0] reducer__in_394;
  wire [15:0] reducer__in_395;
  wire [15:0] reducer__in_396;
  wire [15:0] reducer__in_397;
  wire [15:0] reducer__in_398;
  wire [15:0] reducer__in_399;
  wire [15:0] reducer__in_4;
  wire [15:0] reducer__in_40;
  wire [15:0] reducer__in_400;
  wire [15:0] reducer__in_401;
  wire [15:0] reducer__in_402;
  wire [15:0] reducer__in_403;
  wire [15:0] reducer__in_404;
  wire [15:0] reducer__in_405;
  wire [15:0] reducer__in_406;
  wire [15:0] reducer__in_407;
  wire [15:0] reducer__in_408;
  wire [15:0] reducer__in_409;
  wire [15:0] reducer__in_41;
  wire [15:0] reducer__in_410;
  wire [15:0] reducer__in_411;
  wire [15:0] reducer__in_412;
  wire [15:0] reducer__in_413;
  wire [15:0] reducer__in_414;
  wire [15:0] reducer__in_415;
  wire [15:0] reducer__in_416;
  wire [15:0] reducer__in_417;
  wire [15:0] reducer__in_418;
  wire [15:0] reducer__in_419;
  wire [15:0] reducer__in_42;
  wire [15:0] reducer__in_420;
  wire [15:0] reducer__in_421;
  wire [15:0] reducer__in_422;
  wire [15:0] reducer__in_423;
  wire [15:0] reducer__in_424;
  wire [15:0] reducer__in_425;
  wire [15:0] reducer__in_426;
  wire [15:0] reducer__in_427;
  wire [15:0] reducer__in_428;
  wire [15:0] reducer__in_429;
  wire [15:0] reducer__in_43;
  wire [15:0] reducer__in_430;
  wire [15:0] reducer__in_431;
  wire [15:0] reducer__in_432;
  wire [15:0] reducer__in_433;
  wire [15:0] reducer__in_434;
  wire [15:0] reducer__in_435;
  wire [15:0] reducer__in_436;
  wire [15:0] reducer__in_437;
  wire [15:0] reducer__in_438;
  wire [15:0] reducer__in_439;
  wire [15:0] reducer__in_44;
  wire [15:0] reducer__in_440;
  wire [15:0] reducer__in_441;
  wire [15:0] reducer__in_442;
  wire [15:0] reducer__in_443;
  wire [15:0] reducer__in_444;
  wire [15:0] reducer__in_445;
  wire [15:0] reducer__in_446;
  wire [15:0] reducer__in_447;
  wire [15:0] reducer__in_448;
  wire [15:0] reducer__in_449;
  wire [15:0] reducer__in_45;
  wire [15:0] reducer__in_450;
  wire [15:0] reducer__in_451;
  wire [15:0] reducer__in_452;
  wire [15:0] reducer__in_453;
  wire [15:0] reducer__in_454;
  wire [15:0] reducer__in_455;
  wire [15:0] reducer__in_456;
  wire [15:0] reducer__in_457;
  wire [15:0] reducer__in_458;
  wire [15:0] reducer__in_459;
  wire [15:0] reducer__in_46;
  wire [15:0] reducer__in_460;
  wire [15:0] reducer__in_461;
  wire [15:0] reducer__in_462;
  wire [15:0] reducer__in_463;
  wire [15:0] reducer__in_464;
  wire [15:0] reducer__in_465;
  wire [15:0] reducer__in_466;
  wire [15:0] reducer__in_467;
  wire [15:0] reducer__in_468;
  wire [15:0] reducer__in_469;
  wire [15:0] reducer__in_47;
  wire [15:0] reducer__in_470;
  wire [15:0] reducer__in_471;
  wire [15:0] reducer__in_472;
  wire [15:0] reducer__in_473;
  wire [15:0] reducer__in_474;
  wire [15:0] reducer__in_475;
  wire [15:0] reducer__in_476;
  wire [15:0] reducer__in_477;
  wire [15:0] reducer__in_478;
  wire [15:0] reducer__in_479;
  wire [15:0] reducer__in_48;
  wire [15:0] reducer__in_480;
  wire [15:0] reducer__in_481;
  wire [15:0] reducer__in_482;
  wire [15:0] reducer__in_483;
  wire [15:0] reducer__in_484;
  wire [15:0] reducer__in_485;
  wire [15:0] reducer__in_486;
  wire [15:0] reducer__in_487;
  wire [15:0] reducer__in_488;
  wire [15:0] reducer__in_489;
  wire [15:0] reducer__in_49;
  wire [15:0] reducer__in_490;
  wire [15:0] reducer__in_491;
  wire [15:0] reducer__in_492;
  wire [15:0] reducer__in_493;
  wire [15:0] reducer__in_494;
  wire [15:0] reducer__in_495;
  wire [15:0] reducer__in_496;
  wire [15:0] reducer__in_497;
  wire [15:0] reducer__in_498;
  wire [15:0] reducer__in_499;
  wire [15:0] reducer__in_5;
  wire [15:0] reducer__in_50;
  wire [15:0] reducer__in_500;
  wire [15:0] reducer__in_501;
  wire [15:0] reducer__in_502;
  wire [15:0] reducer__in_503;
  wire [15:0] reducer__in_504;
  wire [15:0] reducer__in_505;
  wire [15:0] reducer__in_506;
  wire [15:0] reducer__in_507;
  wire [15:0] reducer__in_508;
  wire [15:0] reducer__in_509;
  wire [15:0] reducer__in_51;
  wire [15:0] reducer__in_510;
  wire [15:0] reducer__in_511;
  wire [15:0] reducer__in_52;
  wire [15:0] reducer__in_53;
  wire [15:0] reducer__in_54;
  wire [15:0] reducer__in_55;
  wire [15:0] reducer__in_56;
  wire [15:0] reducer__in_57;
  wire [15:0] reducer__in_58;
  wire [15:0] reducer__in_59;
  wire [15:0] reducer__in_6;
  wire [15:0] reducer__in_60;
  wire [15:0] reducer__in_61;
  wire [15:0] reducer__in_62;
  wire [15:0] reducer__in_63;
  wire [15:0] reducer__in_64;
  wire [15:0] reducer__in_65;
  wire [15:0] reducer__in_66;
  wire [15:0] reducer__in_67;
  wire [15:0] reducer__in_68;
  wire [15:0] reducer__in_69;
  wire [15:0] reducer__in_7;
  wire [15:0] reducer__in_70;
  wire [15:0] reducer__in_71;
  wire [15:0] reducer__in_72;
  wire [15:0] reducer__in_73;
  wire [15:0] reducer__in_74;
  wire [15:0] reducer__in_75;
  wire [15:0] reducer__in_76;
  wire [15:0] reducer__in_77;
  wire [15:0] reducer__in_78;
  wire [15:0] reducer__in_79;
  wire [15:0] reducer__in_8;
  wire [15:0] reducer__in_80;
  wire [15:0] reducer__in_81;
  wire [15:0] reducer__in_82;
  wire [15:0] reducer__in_83;
  wire [15:0] reducer__in_84;
  wire [15:0] reducer__in_85;
  wire [15:0] reducer__in_86;
  wire [15:0] reducer__in_87;
  wire [15:0] reducer__in_88;
  wire [15:0] reducer__in_89;
  wire [15:0] reducer__in_9;
  wire [15:0] reducer__in_90;
  wire [15:0] reducer__in_91;
  wire [15:0] reducer__in_92;
  wire [15:0] reducer__in_93;
  wire [15:0] reducer__in_94;
  wire [15:0] reducer__in_95;
  wire [15:0] reducer__in_96;
  wire [15:0] reducer__in_97;
  wire [15:0] reducer__in_98;
  wire [15:0] reducer__in_99;
  wire [15:0] reducer__out;
  reduceParallelPower2Inputs_U2 reducer(
    .in_0(reducer__in_0),
    .in_1(reducer__in_1),
    .in_10(reducer__in_10),
    .in_100(reducer__in_100),
    .in_101(reducer__in_101),
    .in_102(reducer__in_102),
    .in_103(reducer__in_103),
    .in_104(reducer__in_104),
    .in_105(reducer__in_105),
    .in_106(reducer__in_106),
    .in_107(reducer__in_107),
    .in_108(reducer__in_108),
    .in_109(reducer__in_109),
    .in_11(reducer__in_11),
    .in_110(reducer__in_110),
    .in_111(reducer__in_111),
    .in_112(reducer__in_112),
    .in_113(reducer__in_113),
    .in_114(reducer__in_114),
    .in_115(reducer__in_115),
    .in_116(reducer__in_116),
    .in_117(reducer__in_117),
    .in_118(reducer__in_118),
    .in_119(reducer__in_119),
    .in_12(reducer__in_12),
    .in_120(reducer__in_120),
    .in_121(reducer__in_121),
    .in_122(reducer__in_122),
    .in_123(reducer__in_123),
    .in_124(reducer__in_124),
    .in_125(reducer__in_125),
    .in_126(reducer__in_126),
    .in_127(reducer__in_127),
    .in_128(reducer__in_128),
    .in_129(reducer__in_129),
    .in_13(reducer__in_13),
    .in_130(reducer__in_130),
    .in_131(reducer__in_131),
    .in_132(reducer__in_132),
    .in_133(reducer__in_133),
    .in_134(reducer__in_134),
    .in_135(reducer__in_135),
    .in_136(reducer__in_136),
    .in_137(reducer__in_137),
    .in_138(reducer__in_138),
    .in_139(reducer__in_139),
    .in_14(reducer__in_14),
    .in_140(reducer__in_140),
    .in_141(reducer__in_141),
    .in_142(reducer__in_142),
    .in_143(reducer__in_143),
    .in_144(reducer__in_144),
    .in_145(reducer__in_145),
    .in_146(reducer__in_146),
    .in_147(reducer__in_147),
    .in_148(reducer__in_148),
    .in_149(reducer__in_149),
    .in_15(reducer__in_15),
    .in_150(reducer__in_150),
    .in_151(reducer__in_151),
    .in_152(reducer__in_152),
    .in_153(reducer__in_153),
    .in_154(reducer__in_154),
    .in_155(reducer__in_155),
    .in_156(reducer__in_156),
    .in_157(reducer__in_157),
    .in_158(reducer__in_158),
    .in_159(reducer__in_159),
    .in_16(reducer__in_16),
    .in_160(reducer__in_160),
    .in_161(reducer__in_161),
    .in_162(reducer__in_162),
    .in_163(reducer__in_163),
    .in_164(reducer__in_164),
    .in_165(reducer__in_165),
    .in_166(reducer__in_166),
    .in_167(reducer__in_167),
    .in_168(reducer__in_168),
    .in_169(reducer__in_169),
    .in_17(reducer__in_17),
    .in_170(reducer__in_170),
    .in_171(reducer__in_171),
    .in_172(reducer__in_172),
    .in_173(reducer__in_173),
    .in_174(reducer__in_174),
    .in_175(reducer__in_175),
    .in_176(reducer__in_176),
    .in_177(reducer__in_177),
    .in_178(reducer__in_178),
    .in_179(reducer__in_179),
    .in_18(reducer__in_18),
    .in_180(reducer__in_180),
    .in_181(reducer__in_181),
    .in_182(reducer__in_182),
    .in_183(reducer__in_183),
    .in_184(reducer__in_184),
    .in_185(reducer__in_185),
    .in_186(reducer__in_186),
    .in_187(reducer__in_187),
    .in_188(reducer__in_188),
    .in_189(reducer__in_189),
    .in_19(reducer__in_19),
    .in_190(reducer__in_190),
    .in_191(reducer__in_191),
    .in_192(reducer__in_192),
    .in_193(reducer__in_193),
    .in_194(reducer__in_194),
    .in_195(reducer__in_195),
    .in_196(reducer__in_196),
    .in_197(reducer__in_197),
    .in_198(reducer__in_198),
    .in_199(reducer__in_199),
    .in_2(reducer__in_2),
    .in_20(reducer__in_20),
    .in_200(reducer__in_200),
    .in_201(reducer__in_201),
    .in_202(reducer__in_202),
    .in_203(reducer__in_203),
    .in_204(reducer__in_204),
    .in_205(reducer__in_205),
    .in_206(reducer__in_206),
    .in_207(reducer__in_207),
    .in_208(reducer__in_208),
    .in_209(reducer__in_209),
    .in_21(reducer__in_21),
    .in_210(reducer__in_210),
    .in_211(reducer__in_211),
    .in_212(reducer__in_212),
    .in_213(reducer__in_213),
    .in_214(reducer__in_214),
    .in_215(reducer__in_215),
    .in_216(reducer__in_216),
    .in_217(reducer__in_217),
    .in_218(reducer__in_218),
    .in_219(reducer__in_219),
    .in_22(reducer__in_22),
    .in_220(reducer__in_220),
    .in_221(reducer__in_221),
    .in_222(reducer__in_222),
    .in_223(reducer__in_223),
    .in_224(reducer__in_224),
    .in_225(reducer__in_225),
    .in_226(reducer__in_226),
    .in_227(reducer__in_227),
    .in_228(reducer__in_228),
    .in_229(reducer__in_229),
    .in_23(reducer__in_23),
    .in_230(reducer__in_230),
    .in_231(reducer__in_231),
    .in_232(reducer__in_232),
    .in_233(reducer__in_233),
    .in_234(reducer__in_234),
    .in_235(reducer__in_235),
    .in_236(reducer__in_236),
    .in_237(reducer__in_237),
    .in_238(reducer__in_238),
    .in_239(reducer__in_239),
    .in_24(reducer__in_24),
    .in_240(reducer__in_240),
    .in_241(reducer__in_241),
    .in_242(reducer__in_242),
    .in_243(reducer__in_243),
    .in_244(reducer__in_244),
    .in_245(reducer__in_245),
    .in_246(reducer__in_246),
    .in_247(reducer__in_247),
    .in_248(reducer__in_248),
    .in_249(reducer__in_249),
    .in_25(reducer__in_25),
    .in_250(reducer__in_250),
    .in_251(reducer__in_251),
    .in_252(reducer__in_252),
    .in_253(reducer__in_253),
    .in_254(reducer__in_254),
    .in_255(reducer__in_255),
    .in_256(reducer__in_256),
    .in_257(reducer__in_257),
    .in_258(reducer__in_258),
    .in_259(reducer__in_259),
    .in_26(reducer__in_26),
    .in_260(reducer__in_260),
    .in_261(reducer__in_261),
    .in_262(reducer__in_262),
    .in_263(reducer__in_263),
    .in_264(reducer__in_264),
    .in_265(reducer__in_265),
    .in_266(reducer__in_266),
    .in_267(reducer__in_267),
    .in_268(reducer__in_268),
    .in_269(reducer__in_269),
    .in_27(reducer__in_27),
    .in_270(reducer__in_270),
    .in_271(reducer__in_271),
    .in_272(reducer__in_272),
    .in_273(reducer__in_273),
    .in_274(reducer__in_274),
    .in_275(reducer__in_275),
    .in_276(reducer__in_276),
    .in_277(reducer__in_277),
    .in_278(reducer__in_278),
    .in_279(reducer__in_279),
    .in_28(reducer__in_28),
    .in_280(reducer__in_280),
    .in_281(reducer__in_281),
    .in_282(reducer__in_282),
    .in_283(reducer__in_283),
    .in_284(reducer__in_284),
    .in_285(reducer__in_285),
    .in_286(reducer__in_286),
    .in_287(reducer__in_287),
    .in_288(reducer__in_288),
    .in_289(reducer__in_289),
    .in_29(reducer__in_29),
    .in_290(reducer__in_290),
    .in_291(reducer__in_291),
    .in_292(reducer__in_292),
    .in_293(reducer__in_293),
    .in_294(reducer__in_294),
    .in_295(reducer__in_295),
    .in_296(reducer__in_296),
    .in_297(reducer__in_297),
    .in_298(reducer__in_298),
    .in_299(reducer__in_299),
    .in_3(reducer__in_3),
    .in_30(reducer__in_30),
    .in_300(reducer__in_300),
    .in_301(reducer__in_301),
    .in_302(reducer__in_302),
    .in_303(reducer__in_303),
    .in_304(reducer__in_304),
    .in_305(reducer__in_305),
    .in_306(reducer__in_306),
    .in_307(reducer__in_307),
    .in_308(reducer__in_308),
    .in_309(reducer__in_309),
    .in_31(reducer__in_31),
    .in_310(reducer__in_310),
    .in_311(reducer__in_311),
    .in_312(reducer__in_312),
    .in_313(reducer__in_313),
    .in_314(reducer__in_314),
    .in_315(reducer__in_315),
    .in_316(reducer__in_316),
    .in_317(reducer__in_317),
    .in_318(reducer__in_318),
    .in_319(reducer__in_319),
    .in_32(reducer__in_32),
    .in_320(reducer__in_320),
    .in_321(reducer__in_321),
    .in_322(reducer__in_322),
    .in_323(reducer__in_323),
    .in_324(reducer__in_324),
    .in_325(reducer__in_325),
    .in_326(reducer__in_326),
    .in_327(reducer__in_327),
    .in_328(reducer__in_328),
    .in_329(reducer__in_329),
    .in_33(reducer__in_33),
    .in_330(reducer__in_330),
    .in_331(reducer__in_331),
    .in_332(reducer__in_332),
    .in_333(reducer__in_333),
    .in_334(reducer__in_334),
    .in_335(reducer__in_335),
    .in_336(reducer__in_336),
    .in_337(reducer__in_337),
    .in_338(reducer__in_338),
    .in_339(reducer__in_339),
    .in_34(reducer__in_34),
    .in_340(reducer__in_340),
    .in_341(reducer__in_341),
    .in_342(reducer__in_342),
    .in_343(reducer__in_343),
    .in_344(reducer__in_344),
    .in_345(reducer__in_345),
    .in_346(reducer__in_346),
    .in_347(reducer__in_347),
    .in_348(reducer__in_348),
    .in_349(reducer__in_349),
    .in_35(reducer__in_35),
    .in_350(reducer__in_350),
    .in_351(reducer__in_351),
    .in_352(reducer__in_352),
    .in_353(reducer__in_353),
    .in_354(reducer__in_354),
    .in_355(reducer__in_355),
    .in_356(reducer__in_356),
    .in_357(reducer__in_357),
    .in_358(reducer__in_358),
    .in_359(reducer__in_359),
    .in_36(reducer__in_36),
    .in_360(reducer__in_360),
    .in_361(reducer__in_361),
    .in_362(reducer__in_362),
    .in_363(reducer__in_363),
    .in_364(reducer__in_364),
    .in_365(reducer__in_365),
    .in_366(reducer__in_366),
    .in_367(reducer__in_367),
    .in_368(reducer__in_368),
    .in_369(reducer__in_369),
    .in_37(reducer__in_37),
    .in_370(reducer__in_370),
    .in_371(reducer__in_371),
    .in_372(reducer__in_372),
    .in_373(reducer__in_373),
    .in_374(reducer__in_374),
    .in_375(reducer__in_375),
    .in_376(reducer__in_376),
    .in_377(reducer__in_377),
    .in_378(reducer__in_378),
    .in_379(reducer__in_379),
    .in_38(reducer__in_38),
    .in_380(reducer__in_380),
    .in_381(reducer__in_381),
    .in_382(reducer__in_382),
    .in_383(reducer__in_383),
    .in_384(reducer__in_384),
    .in_385(reducer__in_385),
    .in_386(reducer__in_386),
    .in_387(reducer__in_387),
    .in_388(reducer__in_388),
    .in_389(reducer__in_389),
    .in_39(reducer__in_39),
    .in_390(reducer__in_390),
    .in_391(reducer__in_391),
    .in_392(reducer__in_392),
    .in_393(reducer__in_393),
    .in_394(reducer__in_394),
    .in_395(reducer__in_395),
    .in_396(reducer__in_396),
    .in_397(reducer__in_397),
    .in_398(reducer__in_398),
    .in_399(reducer__in_399),
    .in_4(reducer__in_4),
    .in_40(reducer__in_40),
    .in_400(reducer__in_400),
    .in_401(reducer__in_401),
    .in_402(reducer__in_402),
    .in_403(reducer__in_403),
    .in_404(reducer__in_404),
    .in_405(reducer__in_405),
    .in_406(reducer__in_406),
    .in_407(reducer__in_407),
    .in_408(reducer__in_408),
    .in_409(reducer__in_409),
    .in_41(reducer__in_41),
    .in_410(reducer__in_410),
    .in_411(reducer__in_411),
    .in_412(reducer__in_412),
    .in_413(reducer__in_413),
    .in_414(reducer__in_414),
    .in_415(reducer__in_415),
    .in_416(reducer__in_416),
    .in_417(reducer__in_417),
    .in_418(reducer__in_418),
    .in_419(reducer__in_419),
    .in_42(reducer__in_42),
    .in_420(reducer__in_420),
    .in_421(reducer__in_421),
    .in_422(reducer__in_422),
    .in_423(reducer__in_423),
    .in_424(reducer__in_424),
    .in_425(reducer__in_425),
    .in_426(reducer__in_426),
    .in_427(reducer__in_427),
    .in_428(reducer__in_428),
    .in_429(reducer__in_429),
    .in_43(reducer__in_43),
    .in_430(reducer__in_430),
    .in_431(reducer__in_431),
    .in_432(reducer__in_432),
    .in_433(reducer__in_433),
    .in_434(reducer__in_434),
    .in_435(reducer__in_435),
    .in_436(reducer__in_436),
    .in_437(reducer__in_437),
    .in_438(reducer__in_438),
    .in_439(reducer__in_439),
    .in_44(reducer__in_44),
    .in_440(reducer__in_440),
    .in_441(reducer__in_441),
    .in_442(reducer__in_442),
    .in_443(reducer__in_443),
    .in_444(reducer__in_444),
    .in_445(reducer__in_445),
    .in_446(reducer__in_446),
    .in_447(reducer__in_447),
    .in_448(reducer__in_448),
    .in_449(reducer__in_449),
    .in_45(reducer__in_45),
    .in_450(reducer__in_450),
    .in_451(reducer__in_451),
    .in_452(reducer__in_452),
    .in_453(reducer__in_453),
    .in_454(reducer__in_454),
    .in_455(reducer__in_455),
    .in_456(reducer__in_456),
    .in_457(reducer__in_457),
    .in_458(reducer__in_458),
    .in_459(reducer__in_459),
    .in_46(reducer__in_46),
    .in_460(reducer__in_460),
    .in_461(reducer__in_461),
    .in_462(reducer__in_462),
    .in_463(reducer__in_463),
    .in_464(reducer__in_464),
    .in_465(reducer__in_465),
    .in_466(reducer__in_466),
    .in_467(reducer__in_467),
    .in_468(reducer__in_468),
    .in_469(reducer__in_469),
    .in_47(reducer__in_47),
    .in_470(reducer__in_470),
    .in_471(reducer__in_471),
    .in_472(reducer__in_472),
    .in_473(reducer__in_473),
    .in_474(reducer__in_474),
    .in_475(reducer__in_475),
    .in_476(reducer__in_476),
    .in_477(reducer__in_477),
    .in_478(reducer__in_478),
    .in_479(reducer__in_479),
    .in_48(reducer__in_48),
    .in_480(reducer__in_480),
    .in_481(reducer__in_481),
    .in_482(reducer__in_482),
    .in_483(reducer__in_483),
    .in_484(reducer__in_484),
    .in_485(reducer__in_485),
    .in_486(reducer__in_486),
    .in_487(reducer__in_487),
    .in_488(reducer__in_488),
    .in_489(reducer__in_489),
    .in_49(reducer__in_49),
    .in_490(reducer__in_490),
    .in_491(reducer__in_491),
    .in_492(reducer__in_492),
    .in_493(reducer__in_493),
    .in_494(reducer__in_494),
    .in_495(reducer__in_495),
    .in_496(reducer__in_496),
    .in_497(reducer__in_497),
    .in_498(reducer__in_498),
    .in_499(reducer__in_499),
    .in_5(reducer__in_5),
    .in_50(reducer__in_50),
    .in_500(reducer__in_500),
    .in_501(reducer__in_501),
    .in_502(reducer__in_502),
    .in_503(reducer__in_503),
    .in_504(reducer__in_504),
    .in_505(reducer__in_505),
    .in_506(reducer__in_506),
    .in_507(reducer__in_507),
    .in_508(reducer__in_508),
    .in_509(reducer__in_509),
    .in_51(reducer__in_51),
    .in_510(reducer__in_510),
    .in_511(reducer__in_511),
    .in_52(reducer__in_52),
    .in_53(reducer__in_53),
    .in_54(reducer__in_54),
    .in_55(reducer__in_55),
    .in_56(reducer__in_56),
    .in_57(reducer__in_57),
    .in_58(reducer__in_58),
    .in_59(reducer__in_59),
    .in_6(reducer__in_6),
    .in_60(reducer__in_60),
    .in_61(reducer__in_61),
    .in_62(reducer__in_62),
    .in_63(reducer__in_63),
    .in_64(reducer__in_64),
    .in_65(reducer__in_65),
    .in_66(reducer__in_66),
    .in_67(reducer__in_67),
    .in_68(reducer__in_68),
    .in_69(reducer__in_69),
    .in_7(reducer__in_7),
    .in_70(reducer__in_70),
    .in_71(reducer__in_71),
    .in_72(reducer__in_72),
    .in_73(reducer__in_73),
    .in_74(reducer__in_74),
    .in_75(reducer__in_75),
    .in_76(reducer__in_76),
    .in_77(reducer__in_77),
    .in_78(reducer__in_78),
    .in_79(reducer__in_79),
    .in_8(reducer__in_8),
    .in_80(reducer__in_80),
    .in_81(reducer__in_81),
    .in_82(reducer__in_82),
    .in_83(reducer__in_83),
    .in_84(reducer__in_84),
    .in_85(reducer__in_85),
    .in_86(reducer__in_86),
    .in_87(reducer__in_87),
    .in_88(reducer__in_88),
    .in_89(reducer__in_89),
    .in_9(reducer__in_9),
    .in_90(reducer__in_90),
    .in_91(reducer__in_91),
    .in_92(reducer__in_92),
    .in_93(reducer__in_93),
    .in_94(reducer__in_94),
    .in_95(reducer__in_95),
    .in_96(reducer__in_96),
    .in_97(reducer__in_97),
    .in_98(reducer__in_98),
    .in_99(reducer__in_99),
    .out(reducer__out)
  );

  //All the connections
  assign out[15:0] = reducer__out[15:0];
  assign reducer__in_11[15:0] = in_data_11[15:0];
  assign reducer__in_12[15:0] = in_data_12[15:0];
  assign reducer__in_13[15:0] = in_data_13[15:0];
  assign reducer__in_14[15:0] = in_data_14[15:0];
  assign reducer__in_15[15:0] = in_data_15[15:0];
  assign reducer__in_16[15:0] = in_data_16[15:0];
  assign reducer__in_17[15:0] = in_data_17[15:0];
  assign reducer__in_18[15:0] = in_data_18[15:0];
  assign reducer__in_19[15:0] = in_data_19[15:0];
  assign reducer__in_20[15:0] = in_data_20[15:0];
  assign reducer__in_21[15:0] = in_data_21[15:0];
  assign reducer__in_22[15:0] = in_data_22[15:0];
  assign reducer__in_0[15:0] = in_data_0[15:0];
  assign reducer__in_1[15:0] = in_data_1[15:0];
  assign reducer__in_2[15:0] = in_data_2[15:0];
  assign reducer__in_3[15:0] = in_data_3[15:0];
  assign reducer__in_4[15:0] = in_data_4[15:0];
  assign reducer__in_5[15:0] = in_data_5[15:0];
  assign reducer__in_6[15:0] = in_data_6[15:0];
  assign reducer__in_7[15:0] = in_data_7[15:0];
  assign reducer__in_8[15:0] = in_data_8[15:0];
  assign reducer__in_9[15:0] = in_data_9[15:0];
  assign reducer__in_10[15:0] = in_data_10[15:0];
  assign reducer__in_256[15:0] = in_data_256[15:0];
  assign reducer__in_255[15:0] = in_data_255[15:0];
  assign reducer__in_254[15:0] = in_data_254[15:0];
  assign reducer__in_257[15:0] = in_data_257[15:0];
  assign reducer__in_23[15:0] = in_data_23[15:0];
  assign reducer__in_24[15:0] = in_data_24[15:0];
  assign reducer__in_25[15:0] = in_data_25[15:0];
  assign reducer__in_26[15:0] = in_data_26[15:0];
  assign reducer__in_27[15:0] = in_data_27[15:0];
  assign reducer__in_28[15:0] = in_data_28[15:0];
  assign reducer__in_29[15:0] = in_data_29[15:0];
  assign reducer__in_30[15:0] = in_data_30[15:0];
  assign reducer__in_31[15:0] = in_data_31[15:0];
  assign reducer__in_32[15:0] = in_data_32[15:0];
  assign reducer__in_33[15:0] = in_data_33[15:0];
  assign reducer__in_34[15:0] = in_data_34[15:0];
  assign reducer__in_35[15:0] = in_data_35[15:0];
  assign reducer__in_36[15:0] = in_data_36[15:0];
  assign reducer__in_37[15:0] = in_data_37[15:0];
  assign reducer__in_38[15:0] = in_data_38[15:0];
  assign reducer__in_39[15:0] = in_data_39[15:0];
  assign reducer__in_40[15:0] = in_data_40[15:0];
  assign reducer__in_41[15:0] = in_data_41[15:0];
  assign reducer__in_42[15:0] = in_data_42[15:0];
  assign reducer__in_43[15:0] = in_data_43[15:0];
  assign reducer__in_44[15:0] = in_data_44[15:0];
  assign reducer__in_45[15:0] = in_data_45[15:0];
  assign reducer__in_46[15:0] = in_data_46[15:0];
  assign reducer__in_47[15:0] = in_data_47[15:0];
  assign reducer__in_48[15:0] = in_data_48[15:0];
  assign reducer__in_49[15:0] = in_data_49[15:0];
  assign reducer__in_50[15:0] = in_data_50[15:0];
  assign reducer__in_51[15:0] = in_data_51[15:0];
  assign reducer__in_52[15:0] = in_data_52[15:0];
  assign reducer__in_53[15:0] = in_data_53[15:0];
  assign reducer__in_54[15:0] = in_data_54[15:0];
  assign reducer__in_55[15:0] = in_data_55[15:0];
  assign reducer__in_56[15:0] = in_data_56[15:0];
  assign reducer__in_57[15:0] = in_data_57[15:0];
  assign reducer__in_58[15:0] = in_data_58[15:0];
  assign reducer__in_59[15:0] = in_data_59[15:0];
  assign reducer__in_60[15:0] = in_data_60[15:0];
  assign reducer__in_61[15:0] = in_data_61[15:0];
  assign reducer__in_62[15:0] = in_data_62[15:0];
  assign reducer__in_63[15:0] = in_data_63[15:0];
  assign reducer__in_64[15:0] = in_data_64[15:0];
  assign reducer__in_65[15:0] = in_data_65[15:0];
  assign reducer__in_66[15:0] = in_data_66[15:0];
  assign reducer__in_67[15:0] = in_data_67[15:0];
  assign reducer__in_68[15:0] = in_data_68[15:0];
  assign reducer__in_69[15:0] = in_data_69[15:0];
  assign reducer__in_70[15:0] = in_data_70[15:0];
  assign reducer__in_71[15:0] = in_data_71[15:0];
  assign reducer__in_72[15:0] = in_data_72[15:0];
  assign reducer__in_73[15:0] = in_data_73[15:0];
  assign reducer__in_74[15:0] = in_data_74[15:0];
  assign reducer__in_75[15:0] = in_data_75[15:0];
  assign reducer__in_76[15:0] = in_data_76[15:0];
  assign reducer__in_77[15:0] = in_data_77[15:0];
  assign reducer__in_78[15:0] = in_data_78[15:0];
  assign reducer__in_79[15:0] = in_data_79[15:0];
  assign reducer__in_80[15:0] = in_data_80[15:0];
  assign reducer__in_81[15:0] = in_data_81[15:0];
  assign reducer__in_82[15:0] = in_data_82[15:0];
  assign reducer__in_83[15:0] = in_data_83[15:0];
  assign reducer__in_84[15:0] = in_data_84[15:0];
  assign reducer__in_85[15:0] = in_data_85[15:0];
  assign reducer__in_86[15:0] = in_data_86[15:0];
  assign reducer__in_87[15:0] = in_data_87[15:0];
  assign reducer__in_88[15:0] = in_data_88[15:0];
  assign reducer__in_89[15:0] = in_data_89[15:0];
  assign reducer__in_90[15:0] = in_data_90[15:0];
  assign reducer__in_91[15:0] = in_data_91[15:0];
  assign reducer__in_92[15:0] = in_data_92[15:0];
  assign reducer__in_93[15:0] = in_data_93[15:0];
  assign reducer__in_94[15:0] = in_data_94[15:0];
  assign reducer__in_95[15:0] = in_data_95[15:0];
  assign reducer__in_96[15:0] = in_data_96[15:0];
  assign reducer__in_97[15:0] = in_data_97[15:0];
  assign reducer__in_98[15:0] = in_data_98[15:0];
  assign reducer__in_99[15:0] = in_data_99[15:0];
  assign reducer__in_100[15:0] = in_data_100[15:0];
  assign reducer__in_101[15:0] = in_data_101[15:0];
  assign reducer__in_102[15:0] = in_data_102[15:0];
  assign reducer__in_103[15:0] = in_data_103[15:0];
  assign reducer__in_104[15:0] = in_data_104[15:0];
  assign reducer__in_105[15:0] = in_data_105[15:0];
  assign reducer__in_106[15:0] = in_data_106[15:0];
  assign reducer__in_107[15:0] = in_data_107[15:0];
  assign reducer__in_108[15:0] = in_data_108[15:0];
  assign reducer__in_109[15:0] = in_data_109[15:0];
  assign reducer__in_110[15:0] = in_data_110[15:0];
  assign reducer__in_111[15:0] = in_data_111[15:0];
  assign reducer__in_112[15:0] = in_data_112[15:0];
  assign reducer__in_113[15:0] = in_data_113[15:0];
  assign reducer__in_114[15:0] = in_data_114[15:0];
  assign reducer__in_115[15:0] = in_data_115[15:0];
  assign reducer__in_116[15:0] = in_data_116[15:0];
  assign reducer__in_117[15:0] = in_data_117[15:0];
  assign reducer__in_118[15:0] = in_data_118[15:0];
  assign reducer__in_119[15:0] = in_data_119[15:0];
  assign reducer__in_120[15:0] = in_data_120[15:0];
  assign reducer__in_121[15:0] = in_data_121[15:0];
  assign reducer__in_122[15:0] = in_data_122[15:0];
  assign reducer__in_123[15:0] = in_data_123[15:0];
  assign reducer__in_124[15:0] = in_data_124[15:0];
  assign reducer__in_125[15:0] = in_data_125[15:0];
  assign reducer__in_126[15:0] = in_data_126[15:0];
  assign reducer__in_127[15:0] = in_data_127[15:0];
  assign reducer__in_128[15:0] = in_data_128[15:0];
  assign reducer__in_129[15:0] = in_data_129[15:0];
  assign reducer__in_130[15:0] = in_data_130[15:0];
  assign reducer__in_131[15:0] = in_data_131[15:0];
  assign reducer__in_132[15:0] = in_data_132[15:0];
  assign reducer__in_133[15:0] = in_data_133[15:0];
  assign reducer__in_134[15:0] = in_data_134[15:0];
  assign reducer__in_135[15:0] = in_data_135[15:0];
  assign reducer__in_136[15:0] = in_data_136[15:0];
  assign reducer__in_137[15:0] = in_data_137[15:0];
  assign reducer__in_138[15:0] = in_data_138[15:0];
  assign reducer__in_139[15:0] = in_data_139[15:0];
  assign reducer__in_140[15:0] = in_data_140[15:0];
  assign reducer__in_141[15:0] = in_data_141[15:0];
  assign reducer__in_142[15:0] = in_data_142[15:0];
  assign reducer__in_143[15:0] = in_data_143[15:0];
  assign reducer__in_144[15:0] = in_data_144[15:0];
  assign reducer__in_145[15:0] = in_data_145[15:0];
  assign reducer__in_146[15:0] = in_data_146[15:0];
  assign reducer__in_147[15:0] = in_data_147[15:0];
  assign reducer__in_148[15:0] = in_data_148[15:0];
  assign reducer__in_149[15:0] = in_data_149[15:0];
  assign reducer__in_150[15:0] = in_data_150[15:0];
  assign reducer__in_151[15:0] = in_data_151[15:0];
  assign reducer__in_152[15:0] = in_data_152[15:0];
  assign reducer__in_153[15:0] = in_data_153[15:0];
  assign reducer__in_154[15:0] = in_data_154[15:0];
  assign reducer__in_155[15:0] = in_data_155[15:0];
  assign reducer__in_156[15:0] = in_data_156[15:0];
  assign reducer__in_157[15:0] = in_data_157[15:0];
  assign reducer__in_158[15:0] = in_data_158[15:0];
  assign reducer__in_159[15:0] = in_data_159[15:0];
  assign reducer__in_160[15:0] = in_data_160[15:0];
  assign reducer__in_161[15:0] = in_data_161[15:0];
  assign reducer__in_162[15:0] = in_data_162[15:0];
  assign reducer__in_163[15:0] = in_data_163[15:0];
  assign reducer__in_164[15:0] = in_data_164[15:0];
  assign reducer__in_165[15:0] = in_data_165[15:0];
  assign reducer__in_166[15:0] = in_data_166[15:0];
  assign reducer__in_167[15:0] = in_data_167[15:0];
  assign reducer__in_168[15:0] = in_data_168[15:0];
  assign reducer__in_169[15:0] = in_data_169[15:0];
  assign reducer__in_170[15:0] = in_data_170[15:0];
  assign reducer__in_171[15:0] = in_data_171[15:0];
  assign reducer__in_172[15:0] = in_data_172[15:0];
  assign reducer__in_173[15:0] = in_data_173[15:0];
  assign reducer__in_174[15:0] = in_data_174[15:0];
  assign reducer__in_175[15:0] = in_data_175[15:0];
  assign reducer__in_176[15:0] = in_data_176[15:0];
  assign reducer__in_177[15:0] = in_data_177[15:0];
  assign reducer__in_178[15:0] = in_data_178[15:0];
  assign reducer__in_179[15:0] = in_data_179[15:0];
  assign reducer__in_180[15:0] = in_data_180[15:0];
  assign reducer__in_181[15:0] = in_data_181[15:0];
  assign reducer__in_182[15:0] = in_data_182[15:0];
  assign reducer__in_183[15:0] = in_data_183[15:0];
  assign reducer__in_184[15:0] = in_data_184[15:0];
  assign reducer__in_185[15:0] = in_data_185[15:0];
  assign reducer__in_186[15:0] = in_data_186[15:0];
  assign reducer__in_187[15:0] = in_data_187[15:0];
  assign reducer__in_188[15:0] = in_data_188[15:0];
  assign reducer__in_189[15:0] = in_data_189[15:0];
  assign reducer__in_190[15:0] = in_data_190[15:0];
  assign reducer__in_191[15:0] = in_data_191[15:0];
  assign reducer__in_192[15:0] = in_data_192[15:0];
  assign reducer__in_193[15:0] = in_data_193[15:0];
  assign reducer__in_194[15:0] = in_data_194[15:0];
  assign reducer__in_195[15:0] = in_data_195[15:0];
  assign reducer__in_196[15:0] = in_data_196[15:0];
  assign reducer__in_197[15:0] = in_data_197[15:0];
  assign reducer__in_198[15:0] = in_data_198[15:0];
  assign reducer__in_199[15:0] = in_data_199[15:0];
  assign reducer__in_200[15:0] = in_data_200[15:0];
  assign reducer__in_201[15:0] = in_data_201[15:0];
  assign reducer__in_202[15:0] = in_data_202[15:0];
  assign reducer__in_203[15:0] = in_data_203[15:0];
  assign reducer__in_204[15:0] = in_data_204[15:0];
  assign reducer__in_205[15:0] = in_data_205[15:0];
  assign reducer__in_206[15:0] = in_data_206[15:0];
  assign reducer__in_207[15:0] = in_data_207[15:0];
  assign reducer__in_208[15:0] = in_data_208[15:0];
  assign reducer__in_209[15:0] = in_data_209[15:0];
  assign reducer__in_210[15:0] = in_data_210[15:0];
  assign reducer__in_211[15:0] = in_data_211[15:0];
  assign reducer__in_212[15:0] = in_data_212[15:0];
  assign reducer__in_213[15:0] = in_data_213[15:0];
  assign reducer__in_214[15:0] = in_data_214[15:0];
  assign reducer__in_215[15:0] = in_data_215[15:0];
  assign reducer__in_216[15:0] = in_data_216[15:0];
  assign reducer__in_217[15:0] = in_data_217[15:0];
  assign reducer__in_218[15:0] = in_data_218[15:0];
  assign reducer__in_219[15:0] = in_data_219[15:0];
  assign reducer__in_220[15:0] = in_data_220[15:0];
  assign reducer__in_221[15:0] = in_data_221[15:0];
  assign reducer__in_222[15:0] = in_data_222[15:0];
  assign reducer__in_223[15:0] = in_data_223[15:0];
  assign reducer__in_224[15:0] = in_data_224[15:0];
  assign reducer__in_225[15:0] = in_data_225[15:0];
  assign reducer__in_226[15:0] = in_data_226[15:0];
  assign reducer__in_227[15:0] = in_data_227[15:0];
  assign reducer__in_228[15:0] = in_data_228[15:0];
  assign reducer__in_229[15:0] = in_data_229[15:0];
  assign reducer__in_230[15:0] = in_data_230[15:0];
  assign reducer__in_231[15:0] = in_data_231[15:0];
  assign reducer__in_232[15:0] = in_data_232[15:0];
  assign reducer__in_233[15:0] = in_data_233[15:0];
  assign reducer__in_234[15:0] = in_data_234[15:0];
  assign reducer__in_235[15:0] = in_data_235[15:0];
  assign reducer__in_236[15:0] = in_data_236[15:0];
  assign reducer__in_237[15:0] = in_data_237[15:0];
  assign reducer__in_238[15:0] = in_data_238[15:0];
  assign reducer__in_239[15:0] = in_data_239[15:0];
  assign reducer__in_240[15:0] = in_data_240[15:0];
  assign reducer__in_241[15:0] = in_data_241[15:0];
  assign reducer__in_242[15:0] = in_data_242[15:0];
  assign reducer__in_243[15:0] = in_data_243[15:0];
  assign reducer__in_244[15:0] = in_data_244[15:0];
  assign reducer__in_245[15:0] = in_data_245[15:0];
  assign reducer__in_246[15:0] = in_data_246[15:0];
  assign reducer__in_247[15:0] = in_data_247[15:0];
  assign reducer__in_248[15:0] = in_data_248[15:0];
  assign reducer__in_249[15:0] = in_data_249[15:0];
  assign reducer__in_250[15:0] = in_data_250[15:0];
  assign reducer__in_251[15:0] = in_data_251[15:0];
  assign reducer__in_252[15:0] = in_data_252[15:0];
  assign reducer__in_253[15:0] = in_data_253[15:0];
  assign reducer__in_285[15:0] = in_data_285[15:0];
  assign reducer__in_286[15:0] = in_data_286[15:0];
  assign reducer__in_287[15:0] = in_data_287[15:0];
  assign reducer__in_288[15:0] = in_data_288[15:0];
  assign reducer__in_289[15:0] = in_data_289[15:0];
  assign reducer__in_290[15:0] = in_data_290[15:0];
  assign reducer__in_291[15:0] = in_data_291[15:0];
  assign reducer__in_292[15:0] = in_data_292[15:0];
  assign reducer__in_293[15:0] = in_data_293[15:0];
  assign reducer__in_294[15:0] = in_data_294[15:0];
  assign reducer__in_295[15:0] = in_data_295[15:0];
  assign reducer__in_296[15:0] = in_data_296[15:0];
  assign reducer__in_297[15:0] = in_data_297[15:0];
  assign reducer__in_298[15:0] = in_data_298[15:0];
  assign reducer__in_299[15:0] = in_data_299[15:0];
  assign reducer__in_300[15:0] = in_identity[15:0];
  assign reducer__in_301[15:0] = in_identity[15:0];
  assign reducer__in_302[15:0] = in_identity[15:0];
  assign reducer__in_303[15:0] = in_identity[15:0];
  assign reducer__in_304[15:0] = in_identity[15:0];
  assign reducer__in_305[15:0] = in_identity[15:0];
  assign reducer__in_306[15:0] = in_identity[15:0];
  assign reducer__in_307[15:0] = in_identity[15:0];
  assign reducer__in_308[15:0] = in_identity[15:0];
  assign reducer__in_309[15:0] = in_identity[15:0];
  assign reducer__in_310[15:0] = in_identity[15:0];
  assign reducer__in_311[15:0] = in_identity[15:0];
  assign reducer__in_312[15:0] = in_identity[15:0];
  assign reducer__in_313[15:0] = in_identity[15:0];
  assign reducer__in_314[15:0] = in_identity[15:0];
  assign reducer__in_315[15:0] = in_identity[15:0];
  assign reducer__in_316[15:0] = in_identity[15:0];
  assign reducer__in_317[15:0] = in_identity[15:0];
  assign reducer__in_318[15:0] = in_identity[15:0];
  assign reducer__in_319[15:0] = in_identity[15:0];
  assign reducer__in_320[15:0] = in_identity[15:0];
  assign reducer__in_258[15:0] = in_data_258[15:0];
  assign reducer__in_259[15:0] = in_data_259[15:0];
  assign reducer__in_260[15:0] = in_data_260[15:0];
  assign reducer__in_261[15:0] = in_data_261[15:0];
  assign reducer__in_262[15:0] = in_data_262[15:0];
  assign reducer__in_263[15:0] = in_data_263[15:0];
  assign reducer__in_264[15:0] = in_data_264[15:0];
  assign reducer__in_265[15:0] = in_data_265[15:0];
  assign reducer__in_266[15:0] = in_data_266[15:0];
  assign reducer__in_267[15:0] = in_data_267[15:0];
  assign reducer__in_268[15:0] = in_data_268[15:0];
  assign reducer__in_269[15:0] = in_data_269[15:0];
  assign reducer__in_270[15:0] = in_data_270[15:0];
  assign reducer__in_271[15:0] = in_data_271[15:0];
  assign reducer__in_272[15:0] = in_data_272[15:0];
  assign reducer__in_273[15:0] = in_data_273[15:0];
  assign reducer__in_274[15:0] = in_data_274[15:0];
  assign reducer__in_275[15:0] = in_data_275[15:0];
  assign reducer__in_276[15:0] = in_data_276[15:0];
  assign reducer__in_277[15:0] = in_data_277[15:0];
  assign reducer__in_278[15:0] = in_data_278[15:0];
  assign reducer__in_279[15:0] = in_data_279[15:0];
  assign reducer__in_280[15:0] = in_data_280[15:0];
  assign reducer__in_281[15:0] = in_data_281[15:0];
  assign reducer__in_282[15:0] = in_data_282[15:0];
  assign reducer__in_283[15:0] = in_data_283[15:0];
  assign reducer__in_284[15:0] = in_data_284[15:0];
  assign reducer__in_321[15:0] = in_identity[15:0];
  assign reducer__in_322[15:0] = in_identity[15:0];
  assign reducer__in_323[15:0] = in_identity[15:0];
  assign reducer__in_324[15:0] = in_identity[15:0];
  assign reducer__in_325[15:0] = in_identity[15:0];
  assign reducer__in_326[15:0] = in_identity[15:0];
  assign reducer__in_327[15:0] = in_identity[15:0];
  assign reducer__in_328[15:0] = in_identity[15:0];
  assign reducer__in_329[15:0] = in_identity[15:0];
  assign reducer__in_330[15:0] = in_identity[15:0];
  assign reducer__in_331[15:0] = in_identity[15:0];
  assign reducer__in_332[15:0] = in_identity[15:0];
  assign reducer__in_333[15:0] = in_identity[15:0];
  assign reducer__in_334[15:0] = in_identity[15:0];
  assign reducer__in_335[15:0] = in_identity[15:0];
  assign reducer__in_336[15:0] = in_identity[15:0];
  assign reducer__in_337[15:0] = in_identity[15:0];
  assign reducer__in_338[15:0] = in_identity[15:0];
  assign reducer__in_339[15:0] = in_identity[15:0];
  assign reducer__in_340[15:0] = in_identity[15:0];
  assign reducer__in_341[15:0] = in_identity[15:0];
  assign reducer__in_342[15:0] = in_identity[15:0];
  assign reducer__in_343[15:0] = in_identity[15:0];
  assign reducer__in_344[15:0] = in_identity[15:0];
  assign reducer__in_345[15:0] = in_identity[15:0];
  assign reducer__in_346[15:0] = in_identity[15:0];
  assign reducer__in_347[15:0] = in_identity[15:0];
  assign reducer__in_348[15:0] = in_identity[15:0];
  assign reducer__in_349[15:0] = in_identity[15:0];
  assign reducer__in_350[15:0] = in_identity[15:0];
  assign reducer__in_351[15:0] = in_identity[15:0];
  assign reducer__in_352[15:0] = in_identity[15:0];
  assign reducer__in_353[15:0] = in_identity[15:0];
  assign reducer__in_354[15:0] = in_identity[15:0];
  assign reducer__in_355[15:0] = in_identity[15:0];
  assign reducer__in_356[15:0] = in_identity[15:0];
  assign reducer__in_357[15:0] = in_identity[15:0];
  assign reducer__in_358[15:0] = in_identity[15:0];
  assign reducer__in_359[15:0] = in_identity[15:0];
  assign reducer__in_360[15:0] = in_identity[15:0];
  assign reducer__in_361[15:0] = in_identity[15:0];
  assign reducer__in_362[15:0] = in_identity[15:0];
  assign reducer__in_363[15:0] = in_identity[15:0];
  assign reducer__in_364[15:0] = in_identity[15:0];
  assign reducer__in_365[15:0] = in_identity[15:0];
  assign reducer__in_366[15:0] = in_identity[15:0];
  assign reducer__in_367[15:0] = in_identity[15:0];
  assign reducer__in_368[15:0] = in_identity[15:0];
  assign reducer__in_369[15:0] = in_identity[15:0];
  assign reducer__in_370[15:0] = in_identity[15:0];
  assign reducer__in_371[15:0] = in_identity[15:0];
  assign reducer__in_372[15:0] = in_identity[15:0];
  assign reducer__in_373[15:0] = in_identity[15:0];
  assign reducer__in_374[15:0] = in_identity[15:0];
  assign reducer__in_375[15:0] = in_identity[15:0];
  assign reducer__in_376[15:0] = in_identity[15:0];
  assign reducer__in_377[15:0] = in_identity[15:0];
  assign reducer__in_378[15:0] = in_identity[15:0];
  assign reducer__in_379[15:0] = in_identity[15:0];
  assign reducer__in_380[15:0] = in_identity[15:0];
  assign reducer__in_381[15:0] = in_identity[15:0];
  assign reducer__in_382[15:0] = in_identity[15:0];
  assign reducer__in_383[15:0] = in_identity[15:0];
  assign reducer__in_384[15:0] = in_identity[15:0];
  assign reducer__in_385[15:0] = in_identity[15:0];
  assign reducer__in_386[15:0] = in_identity[15:0];
  assign reducer__in_387[15:0] = in_identity[15:0];
  assign reducer__in_388[15:0] = in_identity[15:0];
  assign reducer__in_389[15:0] = in_identity[15:0];
  assign reducer__in_390[15:0] = in_identity[15:0];
  assign reducer__in_391[15:0] = in_identity[15:0];
  assign reducer__in_392[15:0] = in_identity[15:0];
  assign reducer__in_393[15:0] = in_identity[15:0];
  assign reducer__in_394[15:0] = in_identity[15:0];
  assign reducer__in_395[15:0] = in_identity[15:0];
  assign reducer__in_396[15:0] = in_identity[15:0];
  assign reducer__in_397[15:0] = in_identity[15:0];
  assign reducer__in_398[15:0] = in_identity[15:0];
  assign reducer__in_399[15:0] = in_identity[15:0];
  assign reducer__in_400[15:0] = in_identity[15:0];
  assign reducer__in_401[15:0] = in_identity[15:0];
  assign reducer__in_402[15:0] = in_identity[15:0];
  assign reducer__in_403[15:0] = in_identity[15:0];
  assign reducer__in_404[15:0] = in_identity[15:0];
  assign reducer__in_405[15:0] = in_identity[15:0];
  assign reducer__in_406[15:0] = in_identity[15:0];
  assign reducer__in_407[15:0] = in_identity[15:0];
  assign reducer__in_408[15:0] = in_identity[15:0];
  assign reducer__in_409[15:0] = in_identity[15:0];
  assign reducer__in_410[15:0] = in_identity[15:0];
  assign reducer__in_411[15:0] = in_identity[15:0];
  assign reducer__in_412[15:0] = in_identity[15:0];
  assign reducer__in_413[15:0] = in_identity[15:0];
  assign reducer__in_414[15:0] = in_identity[15:0];
  assign reducer__in_415[15:0] = in_identity[15:0];
  assign reducer__in_416[15:0] = in_identity[15:0];
  assign reducer__in_417[15:0] = in_identity[15:0];
  assign reducer__in_418[15:0] = in_identity[15:0];
  assign reducer__in_419[15:0] = in_identity[15:0];
  assign reducer__in_420[15:0] = in_identity[15:0];
  assign reducer__in_421[15:0] = in_identity[15:0];
  assign reducer__in_422[15:0] = in_identity[15:0];
  assign reducer__in_423[15:0] = in_identity[15:0];
  assign reducer__in_424[15:0] = in_identity[15:0];
  assign reducer__in_425[15:0] = in_identity[15:0];
  assign reducer__in_426[15:0] = in_identity[15:0];
  assign reducer__in_427[15:0] = in_identity[15:0];
  assign reducer__in_428[15:0] = in_identity[15:0];
  assign reducer__in_429[15:0] = in_identity[15:0];
  assign reducer__in_430[15:0] = in_identity[15:0];
  assign reducer__in_431[15:0] = in_identity[15:0];
  assign reducer__in_432[15:0] = in_identity[15:0];
  assign reducer__in_433[15:0] = in_identity[15:0];
  assign reducer__in_434[15:0] = in_identity[15:0];
  assign reducer__in_435[15:0] = in_identity[15:0];
  assign reducer__in_436[15:0] = in_identity[15:0];
  assign reducer__in_437[15:0] = in_identity[15:0];
  assign reducer__in_438[15:0] = in_identity[15:0];
  assign reducer__in_439[15:0] = in_identity[15:0];
  assign reducer__in_440[15:0] = in_identity[15:0];
  assign reducer__in_441[15:0] = in_identity[15:0];
  assign reducer__in_442[15:0] = in_identity[15:0];
  assign reducer__in_443[15:0] = in_identity[15:0];
  assign reducer__in_444[15:0] = in_identity[15:0];
  assign reducer__in_445[15:0] = in_identity[15:0];
  assign reducer__in_446[15:0] = in_identity[15:0];
  assign reducer__in_447[15:0] = in_identity[15:0];
  assign reducer__in_448[15:0] = in_identity[15:0];
  assign reducer__in_449[15:0] = in_identity[15:0];
  assign reducer__in_450[15:0] = in_identity[15:0];
  assign reducer__in_451[15:0] = in_identity[15:0];
  assign reducer__in_452[15:0] = in_identity[15:0];
  assign reducer__in_453[15:0] = in_identity[15:0];
  assign reducer__in_454[15:0] = in_identity[15:0];
  assign reducer__in_455[15:0] = in_identity[15:0];
  assign reducer__in_456[15:0] = in_identity[15:0];
  assign reducer__in_457[15:0] = in_identity[15:0];
  assign reducer__in_458[15:0] = in_identity[15:0];
  assign reducer__in_459[15:0] = in_identity[15:0];
  assign reducer__in_460[15:0] = in_identity[15:0];
  assign reducer__in_461[15:0] = in_identity[15:0];
  assign reducer__in_462[15:0] = in_identity[15:0];
  assign reducer__in_463[15:0] = in_identity[15:0];
  assign reducer__in_464[15:0] = in_identity[15:0];
  assign reducer__in_465[15:0] = in_identity[15:0];
  assign reducer__in_466[15:0] = in_identity[15:0];
  assign reducer__in_467[15:0] = in_identity[15:0];
  assign reducer__in_468[15:0] = in_identity[15:0];
  assign reducer__in_469[15:0] = in_identity[15:0];
  assign reducer__in_470[15:0] = in_identity[15:0];
  assign reducer__in_471[15:0] = in_identity[15:0];
  assign reducer__in_472[15:0] = in_identity[15:0];
  assign reducer__in_473[15:0] = in_identity[15:0];
  assign reducer__in_474[15:0] = in_identity[15:0];
  assign reducer__in_475[15:0] = in_identity[15:0];
  assign reducer__in_476[15:0] = in_identity[15:0];
  assign reducer__in_477[15:0] = in_identity[15:0];
  assign reducer__in_478[15:0] = in_identity[15:0];
  assign reducer__in_479[15:0] = in_identity[15:0];
  assign reducer__in_480[15:0] = in_identity[15:0];
  assign reducer__in_481[15:0] = in_identity[15:0];
  assign reducer__in_482[15:0] = in_identity[15:0];
  assign reducer__in_483[15:0] = in_identity[15:0];
  assign reducer__in_484[15:0] = in_identity[15:0];
  assign reducer__in_485[15:0] = in_identity[15:0];
  assign reducer__in_486[15:0] = in_identity[15:0];
  assign reducer__in_487[15:0] = in_identity[15:0];
  assign reducer__in_488[15:0] = in_identity[15:0];
  assign reducer__in_489[15:0] = in_identity[15:0];
  assign reducer__in_490[15:0] = in_identity[15:0];
  assign reducer__in_491[15:0] = in_identity[15:0];
  assign reducer__in_492[15:0] = in_identity[15:0];
  assign reducer__in_493[15:0] = in_identity[15:0];
  assign reducer__in_494[15:0] = in_identity[15:0];
  assign reducer__in_495[15:0] = in_identity[15:0];
  assign reducer__in_496[15:0] = in_identity[15:0];
  assign reducer__in_497[15:0] = in_identity[15:0];
  assign reducer__in_498[15:0] = in_identity[15:0];
  assign reducer__in_499[15:0] = in_identity[15:0];
  assign reducer__in_500[15:0] = in_identity[15:0];
  assign reducer__in_501[15:0] = in_identity[15:0];
  assign reducer__in_502[15:0] = in_identity[15:0];
  assign reducer__in_503[15:0] = in_identity[15:0];
  assign reducer__in_504[15:0] = in_identity[15:0];
  assign reducer__in_505[15:0] = in_identity[15:0];
  assign reducer__in_506[15:0] = in_identity[15:0];
  assign reducer__in_507[15:0] = in_identity[15:0];
  assign reducer__in_508[15:0] = in_identity[15:0];
  assign reducer__in_509[15:0] = in_identity[15:0];
  assign reducer__in_510[15:0] = in_identity[15:0];
  assign reducer__in_511[15:0] = in_identity[15:0];

endmodule //reduceParallel_U1

module reg_U12 #(parameter init=1) (
  input  clk,
  input  clr,
  input  en,
  input [9:0] in,
  output [9:0] out
);
  //Wire declarations for instance 'c0' (Module coreir_const)
  wire [9:0] c0__out;
  coreir_const #(.value(10'b0000000000),.width(10)) c0(
    .out(c0__out)
  );

  //Wire declarations for instance 'clrMux' (Module coreir_mux)
  wire [9:0] clrMux__in0;
  wire [9:0] clrMux__in1;
  wire [9:0] clrMux__out;
  wire  clrMux__sel;
  coreir_mux #(.width(10)) clrMux(
    .in0(clrMux__in0),
    .in1(clrMux__in1),
    .out(clrMux__out),
    .sel(clrMux__sel)
  );

  //Wire declarations for instance 'enMux' (Module coreir_mux)
  wire [9:0] enMux__in0;
  wire [9:0] enMux__in1;
  wire [9:0] enMux__out;
  wire  enMux__sel;
  coreir_mux #(.width(10)) enMux(
    .in0(enMux__in0),
    .in1(enMux__in1),
    .out(enMux__out),
    .sel(enMux__sel)
  );

  //Wire declarations for instance 'reg0' (Module coreir_reg)
  wire  reg0__clk;
  wire [9:0] reg0__in;
  wire [9:0] reg0__out;
  coreir_reg #(.clk_posedge(1),.init(init),.width(10)) reg0(
    .clk(reg0__clk),
    .in(reg0__in),
    .out(reg0__out)
  );

  //All the connections
  assign reg0__in[9:0] = enMux__out[9:0];
  assign out[9:0] = reg0__out[9:0];
  assign enMux__in0[9:0] = reg0__out[9:0];
  assign reg0__clk = clk;
  assign enMux__sel = en;
  assign enMux__in1[9:0] = clrMux__out[9:0];
  assign clrMux__in1[9:0] = c0__out[9:0];
  assign clrMux__sel = clr;
  assign clrMux__in0[9:0] = in[9:0];

endmodule //reg_U12

module reg_U13 #(parameter init=1) (
  input  clk,
  input  clr,
  input  en,
  input [0:0] in,
  output [0:0] out
);
  //Wire declarations for instance 'c0' (Module coreir_const)
  wire [0:0] c0__out;
  coreir_const #(.value(1'b0),.width(1)) c0(
    .out(c0__out)
  );

  //Wire declarations for instance 'clrMux' (Module coreir_mux)
  wire [0:0] clrMux__in0;
  wire [0:0] clrMux__in1;
  wire [0:0] clrMux__out;
  wire  clrMux__sel;
  coreir_mux #(.width(1)) clrMux(
    .in0(clrMux__in0),
    .in1(clrMux__in1),
    .out(clrMux__out),
    .sel(clrMux__sel)
  );

  //Wire declarations for instance 'enMux' (Module coreir_mux)
  wire [0:0] enMux__in0;
  wire [0:0] enMux__in1;
  wire [0:0] enMux__out;
  wire  enMux__sel;
  coreir_mux #(.width(1)) enMux(
    .in0(enMux__in0),
    .in1(enMux__in1),
    .out(enMux__out),
    .sel(enMux__sel)
  );

  //Wire declarations for instance 'reg0' (Module coreir_reg)
  wire  reg0__clk;
  wire [0:0] reg0__in;
  wire [0:0] reg0__out;
  coreir_reg #(.clk_posedge(1),.init(init),.width(1)) reg0(
    .clk(reg0__clk),
    .in(reg0__in),
    .out(reg0__out)
  );

  //All the connections
  assign reg0__in[0:0] = enMux__out[0:0];
  assign out[0:0] = reg0__out[0:0];
  assign enMux__in0[0:0] = reg0__out[0:0];
  assign reg0__clk = clk;
  assign enMux__sel = en;
  assign enMux__in1[0:0] = clrMux__out[0:0];
  assign clrMux__in1[0:0] = c0__out[0:0];
  assign clrMux__sel = clr;
  assign clrMux__in0[0:0] = in[0:0];

endmodule //reg_U13

module rowbuffer_U4 (
  input  clk,
  input  flush,
  output [15:0] rdata,
  output  valid,
  input [15:0] wdata,
  input  wen
);
  //Wire declarations for instance 'add_wen' (Module coreir_add)
  wire [9:0] add_wen__in0;
  wire [9:0] add_wen__in1;
  wire [9:0] add_wen__out;
  coreir_add #(.width(10)) add_wen(
    .in0(add_wen__in0),
    .in1(add_wen__in1),
    .out(add_wen__out)
  );

  //Wire declarations for instance 'c1' (Module corebit_const)
  wire  c1__out;
  corebit_const #(.value(1)) c1(
    .out(c1__out)
  );

  //Wire declarations for instance 'cnt' (Module reg_U12)
  wire  cnt__clk;
  wire  cnt__clr;
  wire  cnt__en;
  wire [9:0] cnt__in;
  wire [9:0] cnt__out;
  reg_U12 #(.init(10'b0000000000)) cnt(
    .clk(cnt__clk),
    .clr(cnt__clr),
    .en(cnt__en),
    .in(cnt__in),
    .out(cnt__out)
  );

  //Wire declarations for instance 'depth_m1' (Module coreir_const)
  wire [9:0] depth_m1__out;
  coreir_const #(.value(10'b0101000000),.width(10)) depth_m1(
    .out(depth_m1__out)
  );

  //Wire declarations for instance 'eq_depth' (Module coreir_eq)
  wire [9:0] eq_depth__in0;
  wire [9:0] eq_depth__in1;
  wire  eq_depth__out;
  coreir_eq #(.width(10)) eq_depth(
    .in0(eq_depth__in0),
    .in1(eq_depth__in1),
    .out(eq_depth__out)
  );

  //Wire declarations for instance 'mem' (Module coreir_mem)
  wire  mem__clk;
  wire [8:0] mem__raddr;
  wire [15:0] mem__rdata;
  wire [8:0] mem__waddr;
  wire [15:0] mem__wdata;
  wire  mem__wen;
  coreir_mem #(.depth(320),.has_init(0),.width(16)) mem(
    .clk(mem__clk),
    .raddr(mem__raddr),
    .rdata(mem__rdata),
    .waddr(mem__waddr),
    .wdata(mem__wdata),
    .wen(mem__wen)
  );

  //Wire declarations for instance 'out_and_wen' (Module corebit_and)
  wire  out_and_wen__in0;
  wire  out_and_wen__in1;
  wire  out_and_wen__out;
  corebit_and out_and_wen(
    .in0(out_and_wen__in0),
    .in1(out_and_wen__in1),
    .out(out_and_wen__out)
  );

  //Wire declarations for instance 'raddr' (Module counter_U11)
  wire  raddr__clk;
  wire  raddr__en;
  wire [8:0] raddr__out;
  wire  raddr__srst;
  counter_U11 #(.init(9'b000000000),.max(9'b100111111)) raddr(
    .clk(raddr__clk),
    .en(raddr__en),
    .out(raddr__out),
    .srst(raddr__srst)
  );

  //Wire declarations for instance 'state' (Module reg_U13)
  wire  state__clk;
  wire  state__clr;
  wire  state__en;
  wire [0:0] state__in;
  wire [0:0] state__out;
  reg_U13 #(.init(1'b0)) state(
    .clk(state__clk),
    .clr(state__clr),
    .en(state__en),
    .in(state__in),
    .out(state__out)
  );

  //Wire declarations for instance 'state0' (Module corebit_not)
  wire  state0__in;
  wire  state0__out;
  corebit_not state0(
    .in(state0__in),
    .out(state0__out)
  );

  //Wire declarations for instance 'waddr' (Module counter_U11)
  wire  waddr__clk;
  wire  waddr__en;
  wire [8:0] waddr__out;
  wire  waddr__srst;
  counter_U11 #(.init(9'b000000000),.max(9'b100111111)) waddr(
    .clk(waddr__clk),
    .en(waddr__en),
    .out(waddr__out),
    .srst(waddr__srst)
  );

  //Wire declarations for instance 'wen_ext' (Module coreir_zext)
  wire [0:0] wen_ext__in;
  wire [9:0] wen_ext__out;
  coreir_zext #(.width_in(1),.width_out(10)) wen_ext(
    .in(wen_ext__in),
    .out(wen_ext__out)
  );

  //All the connections
  assign cnt__clk = clk;
  assign mem__clk = clk;
  assign raddr__clk = clk;
  assign waddr__clk = clk;
  assign state__clk = clk;
  assign mem__raddr[8:0] = raddr__out[8:0];
  assign mem__waddr[8:0] = waddr__out[8:0];
  assign rdata[15:0] = mem__rdata[15:0];
  assign mem__wdata[15:0] = wdata[15:0];
  assign mem__wen = wen;
  assign valid = out_and_wen__out;
  assign raddr__en = out_and_wen__out;
  assign out_and_wen__in1 = wen;
  assign waddr__en = wen;
  assign wen_ext__in[0] = wen;
  assign out_and_wen__in0 = state__out[0];
  assign state0__in = state__out[0];
  assign raddr__srst = flush;
  assign waddr__srst = flush;
  assign cnt__clr = flush;
  assign state__clr = flush;
  assign cnt__en = state0__out;
  assign add_wen__in0[9:0] = wen_ext__out[9:0];
  assign add_wen__in1[9:0] = cnt__out[9:0];
  assign cnt__in[9:0] = add_wen__out[9:0];
  assign eq_depth__in1[9:0] = add_wen__out[9:0];
  assign eq_depth__in0[9:0] = depth_m1__out[9:0];
  assign state__en = eq_depth__out;
  assign state__in[0] = c1__out;

endmodule //rowbuffer_U4

module reg_U20 #(parameter init=1) (
  input  clk,
  input  clr,
  input  en,
  input [15:0] in,
  output [15:0] out
);
  //Wire declarations for instance 'c0' (Module coreir_const)
  wire [15:0] c0__out;
  coreir_const #(.value(16'b0000000000000000),.width(16)) c0(
    .out(c0__out)
  );

  //Wire declarations for instance 'clrMux' (Module coreir_mux)
  wire [15:0] clrMux__in0;
  wire [15:0] clrMux__in1;
  wire [15:0] clrMux__out;
  wire  clrMux__sel;
  coreir_mux #(.width(16)) clrMux(
    .in0(clrMux__in0),
    .in1(clrMux__in1),
    .out(clrMux__out),
    .sel(clrMux__sel)
  );

  //Wire declarations for instance 'enMux' (Module coreir_mux)
  wire [15:0] enMux__in0;
  wire [15:0] enMux__in1;
  wire [15:0] enMux__out;
  wire  enMux__sel;
  coreir_mux #(.width(16)) enMux(
    .in0(enMux__in0),
    .in1(enMux__in1),
    .out(enMux__out),
    .sel(enMux__sel)
  );

  //Wire declarations for instance 'reg0' (Module coreir_reg)
  wire  reg0__clk;
  wire [15:0] reg0__in;
  wire [15:0] reg0__out;
  coreir_reg #(.clk_posedge(1),.init(init),.width(16)) reg0(
    .clk(reg0__clk),
    .in(reg0__in),
    .out(reg0__out)
  );

  //All the connections
  assign reg0__in[15:0] = enMux__out[15:0];
  assign out[15:0] = reg0__out[15:0];
  assign enMux__in0[15:0] = reg0__out[15:0];
  assign reg0__clk = clk;
  assign enMux__sel = en;
  assign enMux__in1[15:0] = clrMux__out[15:0];
  assign clrMux__in1[15:0] = c0__out[15:0];
  assign clrMux__sel = clr;
  assign clrMux__in0[15:0] = in[15:0];

endmodule //reg_U20

module counter_U7 (
  input  clk,
  input  en,
  output [15:0] out,
  output  overflow,
  input  reset
);
  //Wire declarations for instance 'add' (Module coreir_add)
  wire [15:0] add__in0;
  wire [15:0] add__in1;
  wire [15:0] add__out;
  coreir_add #(.width(16)) add(
    .in0(add__in0),
    .in1(add__in1),
    .out(add__out)
  );

  //Wire declarations for instance 'count' (Module reg_U20)
  wire  count__clk;
  wire  count__clr;
  wire  count__en;
  wire [15:0] count__in;
  wire [15:0] count__out;
  reg_U20 #(.init(16'b0000000000000000)) count(
    .clk(count__clk),
    .clr(count__clr),
    .en(count__en),
    .in(count__in),
    .out(count__out)
  );

  //Wire declarations for instance 'inc' (Module coreir_const)
  wire [15:0] inc__out;
  coreir_const #(.value(16'b0000000000000001),.width(16)) inc(
    .out(inc__out)
  );

  //Wire declarations for instance 'max' (Module coreir_const)
  wire [15:0] max__out;
  coreir_const #(.value(16'b0000000100111111),.width(16)) max(
    .out(max__out)
  );

  //Wire declarations for instance 'resetOr' (Module coreir_or)
  wire [0:0] resetOr__in0;
  wire [0:0] resetOr__in1;
  wire [0:0] resetOr__out;
  coreir_or #(.width(1)) resetOr(
    .in0(resetOr__in0),
    .in1(resetOr__in1),
    .out(resetOr__out)
  );

  //Wire declarations for instance 'ult' (Module coreir_ult)
  wire [15:0] ult__in0;
  wire [15:0] ult__in1;
  wire  ult__out;
  coreir_ult #(.width(16)) ult(
    .in0(ult__in0),
    .in1(ult__in1),
    .out(ult__out)
  );

  //All the connections
  assign add__in0[15:0] = count__out[15:0];
  assign out[15:0] = count__out[15:0];
  assign add__in1[15:0] = inc__out[15:0];
  assign count__en = en;
  assign count__in[15:0] = add__out[15:0];
  assign ult__in1[15:0] = add__out[15:0];
  assign ult__in0[15:0] = max__out[15:0];
  assign resetOr__in0[0] = ult__out;
  assign overflow = ult__out;
  assign count__clr = resetOr__out[0];
  assign resetOr__in1[0] = reset;
  assign count__clk = clk;

endmodule //counter_U7

module counter_U8 (
  input  clk,
  input  en,
  output [15:0] out,
  output  overflow,
  input  reset
);
  //Wire declarations for instance 'add' (Module coreir_add)
  wire [15:0] add__in0;
  wire [15:0] add__in1;
  wire [15:0] add__out;
  coreir_add #(.width(16)) add(
    .in0(add__in0),
    .in1(add__in1),
    .out(add__out)
  );

  //Wire declarations for instance 'count' (Module reg_U20)
  wire  count__clk;
  wire  count__clr;
  wire  count__en;
  wire [15:0] count__in;
  wire [15:0] count__out;
  reg_U20 #(.init(16'b0000000000000000)) count(
    .clk(count__clk),
    .clr(count__clr),
    .en(count__en),
    .in(count__in),
    .out(count__out)
  );

  //Wire declarations for instance 'inc' (Module coreir_const)
  wire [15:0] inc__out;
  coreir_const #(.value(16'b0000000000000001),.width(16)) inc(
    .out(inc__out)
  );

  //Wire declarations for instance 'max' (Module coreir_const)
  wire [15:0] max__out;
  coreir_const #(.value(16'b0000000011101111),.width(16)) max(
    .out(max__out)
  );

  //Wire declarations for instance 'resetOr' (Module coreir_or)
  wire [0:0] resetOr__in0;
  wire [0:0] resetOr__in1;
  wire [0:0] resetOr__out;
  coreir_or #(.width(1)) resetOr(
    .in0(resetOr__in0),
    .in1(resetOr__in1),
    .out(resetOr__out)
  );

  //Wire declarations for instance 'ult' (Module coreir_ult)
  wire [15:0] ult__in0;
  wire [15:0] ult__in1;
  wire  ult__out;
  coreir_ult #(.width(16)) ult(
    .in0(ult__in0),
    .in1(ult__in1),
    .out(ult__out)
  );

  //All the connections
  assign add__in0[15:0] = count__out[15:0];
  assign out[15:0] = count__out[15:0];
  assign add__in1[15:0] = inc__out[15:0];
  assign count__en = en;
  assign count__in[15:0] = add__out[15:0];
  assign ult__in1[15:0] = add__out[15:0];
  assign ult__in0[15:0] = max__out[15:0];
  assign resetOr__in0[0] = ult__out;
  assign overflow = ult__out;
  assign count__clr = resetOr__out[0];
  assign resetOr__in1[0] = reset;
  assign count__clk = clk;

endmodule //counter_U8

module linebuffer_U0 (
  input  clk,
  input [15:0] in_0_0,
  output [15:0] out_0_0,
  output [15:0] out_0_1,
  output [15:0] out_0_10,
  output [15:0] out_0_11,
  output [15:0] out_0_12,
  output [15:0] out_0_13,
  output [15:0] out_0_14,
  output [15:0] out_0_15,
  output [15:0] out_0_16,
  output [15:0] out_0_17,
  output [15:0] out_0_18,
  output [15:0] out_0_19,
  output [15:0] out_0_2,
  output [15:0] out_0_3,
  output [15:0] out_0_4,
  output [15:0] out_0_5,
  output [15:0] out_0_6,
  output [15:0] out_0_7,
  output [15:0] out_0_8,
  output [15:0] out_0_9,
  output [15:0] out_10_0,
  output [15:0] out_10_1,
  output [15:0] out_10_10,
  output [15:0] out_10_11,
  output [15:0] out_10_12,
  output [15:0] out_10_13,
  output [15:0] out_10_14,
  output [15:0] out_10_15,
  output [15:0] out_10_16,
  output [15:0] out_10_17,
  output [15:0] out_10_18,
  output [15:0] out_10_19,
  output [15:0] out_10_2,
  output [15:0] out_10_3,
  output [15:0] out_10_4,
  output [15:0] out_10_5,
  output [15:0] out_10_6,
  output [15:0] out_10_7,
  output [15:0] out_10_8,
  output [15:0] out_10_9,
  output [15:0] out_11_0,
  output [15:0] out_11_1,
  output [15:0] out_11_10,
  output [15:0] out_11_11,
  output [15:0] out_11_12,
  output [15:0] out_11_13,
  output [15:0] out_11_14,
  output [15:0] out_11_15,
  output [15:0] out_11_16,
  output [15:0] out_11_17,
  output [15:0] out_11_18,
  output [15:0] out_11_19,
  output [15:0] out_11_2,
  output [15:0] out_11_3,
  output [15:0] out_11_4,
  output [15:0] out_11_5,
  output [15:0] out_11_6,
  output [15:0] out_11_7,
  output [15:0] out_11_8,
  output [15:0] out_11_9,
  output [15:0] out_12_0,
  output [15:0] out_12_1,
  output [15:0] out_12_10,
  output [15:0] out_12_11,
  output [15:0] out_12_12,
  output [15:0] out_12_13,
  output [15:0] out_12_14,
  output [15:0] out_12_15,
  output [15:0] out_12_16,
  output [15:0] out_12_17,
  output [15:0] out_12_18,
  output [15:0] out_12_19,
  output [15:0] out_12_2,
  output [15:0] out_12_3,
  output [15:0] out_12_4,
  output [15:0] out_12_5,
  output [15:0] out_12_6,
  output [15:0] out_12_7,
  output [15:0] out_12_8,
  output [15:0] out_12_9,
  output [15:0] out_13_0,
  output [15:0] out_13_1,
  output [15:0] out_13_10,
  output [15:0] out_13_11,
  output [15:0] out_13_12,
  output [15:0] out_13_13,
  output [15:0] out_13_14,
  output [15:0] out_13_15,
  output [15:0] out_13_16,
  output [15:0] out_13_17,
  output [15:0] out_13_18,
  output [15:0] out_13_19,
  output [15:0] out_13_2,
  output [15:0] out_13_3,
  output [15:0] out_13_4,
  output [15:0] out_13_5,
  output [15:0] out_13_6,
  output [15:0] out_13_7,
  output [15:0] out_13_8,
  output [15:0] out_13_9,
  output [15:0] out_14_0,
  output [15:0] out_14_1,
  output [15:0] out_14_10,
  output [15:0] out_14_11,
  output [15:0] out_14_12,
  output [15:0] out_14_13,
  output [15:0] out_14_14,
  output [15:0] out_14_15,
  output [15:0] out_14_16,
  output [15:0] out_14_17,
  output [15:0] out_14_18,
  output [15:0] out_14_19,
  output [15:0] out_14_2,
  output [15:0] out_14_3,
  output [15:0] out_14_4,
  output [15:0] out_14_5,
  output [15:0] out_14_6,
  output [15:0] out_14_7,
  output [15:0] out_14_8,
  output [15:0] out_14_9,
  output [15:0] out_15_0,
  output [15:0] out_15_1,
  output [15:0] out_15_10,
  output [15:0] out_15_11,
  output [15:0] out_15_12,
  output [15:0] out_15_13,
  output [15:0] out_15_14,
  output [15:0] out_15_15,
  output [15:0] out_15_16,
  output [15:0] out_15_17,
  output [15:0] out_15_18,
  output [15:0] out_15_19,
  output [15:0] out_15_2,
  output [15:0] out_15_3,
  output [15:0] out_15_4,
  output [15:0] out_15_5,
  output [15:0] out_15_6,
  output [15:0] out_15_7,
  output [15:0] out_15_8,
  output [15:0] out_15_9,
  output [15:0] out_1_0,
  output [15:0] out_1_1,
  output [15:0] out_1_10,
  output [15:0] out_1_11,
  output [15:0] out_1_12,
  output [15:0] out_1_13,
  output [15:0] out_1_14,
  output [15:0] out_1_15,
  output [15:0] out_1_16,
  output [15:0] out_1_17,
  output [15:0] out_1_18,
  output [15:0] out_1_19,
  output [15:0] out_1_2,
  output [15:0] out_1_3,
  output [15:0] out_1_4,
  output [15:0] out_1_5,
  output [15:0] out_1_6,
  output [15:0] out_1_7,
  output [15:0] out_1_8,
  output [15:0] out_1_9,
  output [15:0] out_2_0,
  output [15:0] out_2_1,
  output [15:0] out_2_10,
  output [15:0] out_2_11,
  output [15:0] out_2_12,
  output [15:0] out_2_13,
  output [15:0] out_2_14,
  output [15:0] out_2_15,
  output [15:0] out_2_16,
  output [15:0] out_2_17,
  output [15:0] out_2_18,
  output [15:0] out_2_19,
  output [15:0] out_2_2,
  output [15:0] out_2_3,
  output [15:0] out_2_4,
  output [15:0] out_2_5,
  output [15:0] out_2_6,
  output [15:0] out_2_7,
  output [15:0] out_2_8,
  output [15:0] out_2_9,
  output [15:0] out_3_0,
  output [15:0] out_3_1,
  output [15:0] out_3_10,
  output [15:0] out_3_11,
  output [15:0] out_3_12,
  output [15:0] out_3_13,
  output [15:0] out_3_14,
  output [15:0] out_3_15,
  output [15:0] out_3_16,
  output [15:0] out_3_17,
  output [15:0] out_3_18,
  output [15:0] out_3_19,
  output [15:0] out_3_2,
  output [15:0] out_3_3,
  output [15:0] out_3_4,
  output [15:0] out_3_5,
  output [15:0] out_3_6,
  output [15:0] out_3_7,
  output [15:0] out_3_8,
  output [15:0] out_3_9,
  output [15:0] out_4_0,
  output [15:0] out_4_1,
  output [15:0] out_4_10,
  output [15:0] out_4_11,
  output [15:0] out_4_12,
  output [15:0] out_4_13,
  output [15:0] out_4_14,
  output [15:0] out_4_15,
  output [15:0] out_4_16,
  output [15:0] out_4_17,
  output [15:0] out_4_18,
  output [15:0] out_4_19,
  output [15:0] out_4_2,
  output [15:0] out_4_3,
  output [15:0] out_4_4,
  output [15:0] out_4_5,
  output [15:0] out_4_6,
  output [15:0] out_4_7,
  output [15:0] out_4_8,
  output [15:0] out_4_9,
  output [15:0] out_5_0,
  output [15:0] out_5_1,
  output [15:0] out_5_10,
  output [15:0] out_5_11,
  output [15:0] out_5_12,
  output [15:0] out_5_13,
  output [15:0] out_5_14,
  output [15:0] out_5_15,
  output [15:0] out_5_16,
  output [15:0] out_5_17,
  output [15:0] out_5_18,
  output [15:0] out_5_19,
  output [15:0] out_5_2,
  output [15:0] out_5_3,
  output [15:0] out_5_4,
  output [15:0] out_5_5,
  output [15:0] out_5_6,
  output [15:0] out_5_7,
  output [15:0] out_5_8,
  output [15:0] out_5_9,
  output [15:0] out_6_0,
  output [15:0] out_6_1,
  output [15:0] out_6_10,
  output [15:0] out_6_11,
  output [15:0] out_6_12,
  output [15:0] out_6_13,
  output [15:0] out_6_14,
  output [15:0] out_6_15,
  output [15:0] out_6_16,
  output [15:0] out_6_17,
  output [15:0] out_6_18,
  output [15:0] out_6_19,
  output [15:0] out_6_2,
  output [15:0] out_6_3,
  output [15:0] out_6_4,
  output [15:0] out_6_5,
  output [15:0] out_6_6,
  output [15:0] out_6_7,
  output [15:0] out_6_8,
  output [15:0] out_6_9,
  output [15:0] out_7_0,
  output [15:0] out_7_1,
  output [15:0] out_7_10,
  output [15:0] out_7_11,
  output [15:0] out_7_12,
  output [15:0] out_7_13,
  output [15:0] out_7_14,
  output [15:0] out_7_15,
  output [15:0] out_7_16,
  output [15:0] out_7_17,
  output [15:0] out_7_18,
  output [15:0] out_7_19,
  output [15:0] out_7_2,
  output [15:0] out_7_3,
  output [15:0] out_7_4,
  output [15:0] out_7_5,
  output [15:0] out_7_6,
  output [15:0] out_7_7,
  output [15:0] out_7_8,
  output [15:0] out_7_9,
  output [15:0] out_8_0,
  output [15:0] out_8_1,
  output [15:0] out_8_10,
  output [15:0] out_8_11,
  output [15:0] out_8_12,
  output [15:0] out_8_13,
  output [15:0] out_8_14,
  output [15:0] out_8_15,
  output [15:0] out_8_16,
  output [15:0] out_8_17,
  output [15:0] out_8_18,
  output [15:0] out_8_19,
  output [15:0] out_8_2,
  output [15:0] out_8_3,
  output [15:0] out_8_4,
  output [15:0] out_8_5,
  output [15:0] out_8_6,
  output [15:0] out_8_7,
  output [15:0] out_8_8,
  output [15:0] out_8_9,
  output [15:0] out_9_0,
  output [15:0] out_9_1,
  output [15:0] out_9_10,
  output [15:0] out_9_11,
  output [15:0] out_9_12,
  output [15:0] out_9_13,
  output [15:0] out_9_14,
  output [15:0] out_9_15,
  output [15:0] out_9_16,
  output [15:0] out_9_17,
  output [15:0] out_9_18,
  output [15:0] out_9_19,
  output [15:0] out_9_2,
  output [15:0] out_9_3,
  output [15:0] out_9_4,
  output [15:0] out_9_5,
  output [15:0] out_9_6,
  output [15:0] out_9_7,
  output [15:0] out_9_8,
  output [15:0] out_9_9,
  output  valid,
  output  valid_chain,
  input  wen
);
  //Wire declarations for instance 'const_stencil0' (Module coreir_const)
  wire [15:0] const_stencil0__out;
  coreir_const #(.value(16'b0000000000010011),.width(16)) const_stencil0(
    .out(const_stencil0__out)
  );

  //Wire declarations for instance 'const_stencil1' (Module coreir_const)
  wire [15:0] const_stencil1__out;
  coreir_const #(.value(16'b0000000000001111),.width(16)) const_stencil1(
    .out(const_stencil1__out)
  );

  //Wire declarations for instance 'lb1d_0' (Module linebuffer_U3)
  wire  lb1d_0__clk;
  wire [15:0] lb1d_0__in_0;
  wire [15:0] lb1d_0__out_0;
  wire [15:0] lb1d_0__out_1;
  wire [15:0] lb1d_0__out_10;
  wire [15:0] lb1d_0__out_11;
  wire [15:0] lb1d_0__out_12;
  wire [15:0] lb1d_0__out_13;
  wire [15:0] lb1d_0__out_14;
  wire [15:0] lb1d_0__out_15;
  wire [15:0] lb1d_0__out_16;
  wire [15:0] lb1d_0__out_17;
  wire [15:0] lb1d_0__out_18;
  wire [15:0] lb1d_0__out_19;
  wire [15:0] lb1d_0__out_2;
  wire [15:0] lb1d_0__out_3;
  wire [15:0] lb1d_0__out_4;
  wire [15:0] lb1d_0__out_5;
  wire [15:0] lb1d_0__out_6;
  wire [15:0] lb1d_0__out_7;
  wire [15:0] lb1d_0__out_8;
  wire [15:0] lb1d_0__out_9;
  wire  lb1d_0__valid;
  wire  lb1d_0__valid_chain;
  wire  lb1d_0__wen;
  linebuffer_U3 lb1d_0(
    .clk(lb1d_0__clk),
    .in_0(lb1d_0__in_0),
    .out_0(lb1d_0__out_0),
    .out_1(lb1d_0__out_1),
    .out_10(lb1d_0__out_10),
    .out_11(lb1d_0__out_11),
    .out_12(lb1d_0__out_12),
    .out_13(lb1d_0__out_13),
    .out_14(lb1d_0__out_14),
    .out_15(lb1d_0__out_15),
    .out_16(lb1d_0__out_16),
    .out_17(lb1d_0__out_17),
    .out_18(lb1d_0__out_18),
    .out_19(lb1d_0__out_19),
    .out_2(lb1d_0__out_2),
    .out_3(lb1d_0__out_3),
    .out_4(lb1d_0__out_4),
    .out_5(lb1d_0__out_5),
    .out_6(lb1d_0__out_6),
    .out_7(lb1d_0__out_7),
    .out_8(lb1d_0__out_8),
    .out_9(lb1d_0__out_9),
    .valid(lb1d_0__valid),
    .valid_chain(lb1d_0__valid_chain),
    .wen(lb1d_0__wen)
  );

  //Wire declarations for instance 'lb1d_1' (Module linebuffer_U3)
  wire  lb1d_1__clk;
  wire [15:0] lb1d_1__in_0;
  wire [15:0] lb1d_1__out_0;
  wire [15:0] lb1d_1__out_1;
  wire [15:0] lb1d_1__out_10;
  wire [15:0] lb1d_1__out_11;
  wire [15:0] lb1d_1__out_12;
  wire [15:0] lb1d_1__out_13;
  wire [15:0] lb1d_1__out_14;
  wire [15:0] lb1d_1__out_15;
  wire [15:0] lb1d_1__out_16;
  wire [15:0] lb1d_1__out_17;
  wire [15:0] lb1d_1__out_18;
  wire [15:0] lb1d_1__out_19;
  wire [15:0] lb1d_1__out_2;
  wire [15:0] lb1d_1__out_3;
  wire [15:0] lb1d_1__out_4;
  wire [15:0] lb1d_1__out_5;
  wire [15:0] lb1d_1__out_6;
  wire [15:0] lb1d_1__out_7;
  wire [15:0] lb1d_1__out_8;
  wire [15:0] lb1d_1__out_9;
  wire  lb1d_1__valid;
  wire  lb1d_1__valid_chain;
  wire  lb1d_1__wen;
  linebuffer_U3 lb1d_1(
    .clk(lb1d_1__clk),
    .in_0(lb1d_1__in_0),
    .out_0(lb1d_1__out_0),
    .out_1(lb1d_1__out_1),
    .out_10(lb1d_1__out_10),
    .out_11(lb1d_1__out_11),
    .out_12(lb1d_1__out_12),
    .out_13(lb1d_1__out_13),
    .out_14(lb1d_1__out_14),
    .out_15(lb1d_1__out_15),
    .out_16(lb1d_1__out_16),
    .out_17(lb1d_1__out_17),
    .out_18(lb1d_1__out_18),
    .out_19(lb1d_1__out_19),
    .out_2(lb1d_1__out_2),
    .out_3(lb1d_1__out_3),
    .out_4(lb1d_1__out_4),
    .out_5(lb1d_1__out_5),
    .out_6(lb1d_1__out_6),
    .out_7(lb1d_1__out_7),
    .out_8(lb1d_1__out_8),
    .out_9(lb1d_1__out_9),
    .valid(lb1d_1__valid),
    .valid_chain(lb1d_1__valid_chain),
    .wen(lb1d_1__wen)
  );

  //Wire declarations for instance 'lb1d_10' (Module linebuffer_U3)
  wire  lb1d_10__clk;
  wire [15:0] lb1d_10__in_0;
  wire [15:0] lb1d_10__out_0;
  wire [15:0] lb1d_10__out_1;
  wire [15:0] lb1d_10__out_10;
  wire [15:0] lb1d_10__out_11;
  wire [15:0] lb1d_10__out_12;
  wire [15:0] lb1d_10__out_13;
  wire [15:0] lb1d_10__out_14;
  wire [15:0] lb1d_10__out_15;
  wire [15:0] lb1d_10__out_16;
  wire [15:0] lb1d_10__out_17;
  wire [15:0] lb1d_10__out_18;
  wire [15:0] lb1d_10__out_19;
  wire [15:0] lb1d_10__out_2;
  wire [15:0] lb1d_10__out_3;
  wire [15:0] lb1d_10__out_4;
  wire [15:0] lb1d_10__out_5;
  wire [15:0] lb1d_10__out_6;
  wire [15:0] lb1d_10__out_7;
  wire [15:0] lb1d_10__out_8;
  wire [15:0] lb1d_10__out_9;
  wire  lb1d_10__valid;
  wire  lb1d_10__valid_chain;
  wire  lb1d_10__wen;
  linebuffer_U3 lb1d_10(
    .clk(lb1d_10__clk),
    .in_0(lb1d_10__in_0),
    .out_0(lb1d_10__out_0),
    .out_1(lb1d_10__out_1),
    .out_10(lb1d_10__out_10),
    .out_11(lb1d_10__out_11),
    .out_12(lb1d_10__out_12),
    .out_13(lb1d_10__out_13),
    .out_14(lb1d_10__out_14),
    .out_15(lb1d_10__out_15),
    .out_16(lb1d_10__out_16),
    .out_17(lb1d_10__out_17),
    .out_18(lb1d_10__out_18),
    .out_19(lb1d_10__out_19),
    .out_2(lb1d_10__out_2),
    .out_3(lb1d_10__out_3),
    .out_4(lb1d_10__out_4),
    .out_5(lb1d_10__out_5),
    .out_6(lb1d_10__out_6),
    .out_7(lb1d_10__out_7),
    .out_8(lb1d_10__out_8),
    .out_9(lb1d_10__out_9),
    .valid(lb1d_10__valid),
    .valid_chain(lb1d_10__valid_chain),
    .wen(lb1d_10__wen)
  );

  //Wire declarations for instance 'lb1d_11' (Module linebuffer_U3)
  wire  lb1d_11__clk;
  wire [15:0] lb1d_11__in_0;
  wire [15:0] lb1d_11__out_0;
  wire [15:0] lb1d_11__out_1;
  wire [15:0] lb1d_11__out_10;
  wire [15:0] lb1d_11__out_11;
  wire [15:0] lb1d_11__out_12;
  wire [15:0] lb1d_11__out_13;
  wire [15:0] lb1d_11__out_14;
  wire [15:0] lb1d_11__out_15;
  wire [15:0] lb1d_11__out_16;
  wire [15:0] lb1d_11__out_17;
  wire [15:0] lb1d_11__out_18;
  wire [15:0] lb1d_11__out_19;
  wire [15:0] lb1d_11__out_2;
  wire [15:0] lb1d_11__out_3;
  wire [15:0] lb1d_11__out_4;
  wire [15:0] lb1d_11__out_5;
  wire [15:0] lb1d_11__out_6;
  wire [15:0] lb1d_11__out_7;
  wire [15:0] lb1d_11__out_8;
  wire [15:0] lb1d_11__out_9;
  wire  lb1d_11__valid;
  wire  lb1d_11__valid_chain;
  wire  lb1d_11__wen;
  linebuffer_U3 lb1d_11(
    .clk(lb1d_11__clk),
    .in_0(lb1d_11__in_0),
    .out_0(lb1d_11__out_0),
    .out_1(lb1d_11__out_1),
    .out_10(lb1d_11__out_10),
    .out_11(lb1d_11__out_11),
    .out_12(lb1d_11__out_12),
    .out_13(lb1d_11__out_13),
    .out_14(lb1d_11__out_14),
    .out_15(lb1d_11__out_15),
    .out_16(lb1d_11__out_16),
    .out_17(lb1d_11__out_17),
    .out_18(lb1d_11__out_18),
    .out_19(lb1d_11__out_19),
    .out_2(lb1d_11__out_2),
    .out_3(lb1d_11__out_3),
    .out_4(lb1d_11__out_4),
    .out_5(lb1d_11__out_5),
    .out_6(lb1d_11__out_6),
    .out_7(lb1d_11__out_7),
    .out_8(lb1d_11__out_8),
    .out_9(lb1d_11__out_9),
    .valid(lb1d_11__valid),
    .valid_chain(lb1d_11__valid_chain),
    .wen(lb1d_11__wen)
  );

  //Wire declarations for instance 'lb1d_12' (Module linebuffer_U3)
  wire  lb1d_12__clk;
  wire [15:0] lb1d_12__in_0;
  wire [15:0] lb1d_12__out_0;
  wire [15:0] lb1d_12__out_1;
  wire [15:0] lb1d_12__out_10;
  wire [15:0] lb1d_12__out_11;
  wire [15:0] lb1d_12__out_12;
  wire [15:0] lb1d_12__out_13;
  wire [15:0] lb1d_12__out_14;
  wire [15:0] lb1d_12__out_15;
  wire [15:0] lb1d_12__out_16;
  wire [15:0] lb1d_12__out_17;
  wire [15:0] lb1d_12__out_18;
  wire [15:0] lb1d_12__out_19;
  wire [15:0] lb1d_12__out_2;
  wire [15:0] lb1d_12__out_3;
  wire [15:0] lb1d_12__out_4;
  wire [15:0] lb1d_12__out_5;
  wire [15:0] lb1d_12__out_6;
  wire [15:0] lb1d_12__out_7;
  wire [15:0] lb1d_12__out_8;
  wire [15:0] lb1d_12__out_9;
  wire  lb1d_12__valid;
  wire  lb1d_12__valid_chain;
  wire  lb1d_12__wen;
  linebuffer_U3 lb1d_12(
    .clk(lb1d_12__clk),
    .in_0(lb1d_12__in_0),
    .out_0(lb1d_12__out_0),
    .out_1(lb1d_12__out_1),
    .out_10(lb1d_12__out_10),
    .out_11(lb1d_12__out_11),
    .out_12(lb1d_12__out_12),
    .out_13(lb1d_12__out_13),
    .out_14(lb1d_12__out_14),
    .out_15(lb1d_12__out_15),
    .out_16(lb1d_12__out_16),
    .out_17(lb1d_12__out_17),
    .out_18(lb1d_12__out_18),
    .out_19(lb1d_12__out_19),
    .out_2(lb1d_12__out_2),
    .out_3(lb1d_12__out_3),
    .out_4(lb1d_12__out_4),
    .out_5(lb1d_12__out_5),
    .out_6(lb1d_12__out_6),
    .out_7(lb1d_12__out_7),
    .out_8(lb1d_12__out_8),
    .out_9(lb1d_12__out_9),
    .valid(lb1d_12__valid),
    .valid_chain(lb1d_12__valid_chain),
    .wen(lb1d_12__wen)
  );

  //Wire declarations for instance 'lb1d_13' (Module linebuffer_U3)
  wire  lb1d_13__clk;
  wire [15:0] lb1d_13__in_0;
  wire [15:0] lb1d_13__out_0;
  wire [15:0] lb1d_13__out_1;
  wire [15:0] lb1d_13__out_10;
  wire [15:0] lb1d_13__out_11;
  wire [15:0] lb1d_13__out_12;
  wire [15:0] lb1d_13__out_13;
  wire [15:0] lb1d_13__out_14;
  wire [15:0] lb1d_13__out_15;
  wire [15:0] lb1d_13__out_16;
  wire [15:0] lb1d_13__out_17;
  wire [15:0] lb1d_13__out_18;
  wire [15:0] lb1d_13__out_19;
  wire [15:0] lb1d_13__out_2;
  wire [15:0] lb1d_13__out_3;
  wire [15:0] lb1d_13__out_4;
  wire [15:0] lb1d_13__out_5;
  wire [15:0] lb1d_13__out_6;
  wire [15:0] lb1d_13__out_7;
  wire [15:0] lb1d_13__out_8;
  wire [15:0] lb1d_13__out_9;
  wire  lb1d_13__valid;
  wire  lb1d_13__valid_chain;
  wire  lb1d_13__wen;
  linebuffer_U3 lb1d_13(
    .clk(lb1d_13__clk),
    .in_0(lb1d_13__in_0),
    .out_0(lb1d_13__out_0),
    .out_1(lb1d_13__out_1),
    .out_10(lb1d_13__out_10),
    .out_11(lb1d_13__out_11),
    .out_12(lb1d_13__out_12),
    .out_13(lb1d_13__out_13),
    .out_14(lb1d_13__out_14),
    .out_15(lb1d_13__out_15),
    .out_16(lb1d_13__out_16),
    .out_17(lb1d_13__out_17),
    .out_18(lb1d_13__out_18),
    .out_19(lb1d_13__out_19),
    .out_2(lb1d_13__out_2),
    .out_3(lb1d_13__out_3),
    .out_4(lb1d_13__out_4),
    .out_5(lb1d_13__out_5),
    .out_6(lb1d_13__out_6),
    .out_7(lb1d_13__out_7),
    .out_8(lb1d_13__out_8),
    .out_9(lb1d_13__out_9),
    .valid(lb1d_13__valid),
    .valid_chain(lb1d_13__valid_chain),
    .wen(lb1d_13__wen)
  );

  //Wire declarations for instance 'lb1d_14' (Module linebuffer_U3)
  wire  lb1d_14__clk;
  wire [15:0] lb1d_14__in_0;
  wire [15:0] lb1d_14__out_0;
  wire [15:0] lb1d_14__out_1;
  wire [15:0] lb1d_14__out_10;
  wire [15:0] lb1d_14__out_11;
  wire [15:0] lb1d_14__out_12;
  wire [15:0] lb1d_14__out_13;
  wire [15:0] lb1d_14__out_14;
  wire [15:0] lb1d_14__out_15;
  wire [15:0] lb1d_14__out_16;
  wire [15:0] lb1d_14__out_17;
  wire [15:0] lb1d_14__out_18;
  wire [15:0] lb1d_14__out_19;
  wire [15:0] lb1d_14__out_2;
  wire [15:0] lb1d_14__out_3;
  wire [15:0] lb1d_14__out_4;
  wire [15:0] lb1d_14__out_5;
  wire [15:0] lb1d_14__out_6;
  wire [15:0] lb1d_14__out_7;
  wire [15:0] lb1d_14__out_8;
  wire [15:0] lb1d_14__out_9;
  wire  lb1d_14__valid;
  wire  lb1d_14__valid_chain;
  wire  lb1d_14__wen;
  linebuffer_U3 lb1d_14(
    .clk(lb1d_14__clk),
    .in_0(lb1d_14__in_0),
    .out_0(lb1d_14__out_0),
    .out_1(lb1d_14__out_1),
    .out_10(lb1d_14__out_10),
    .out_11(lb1d_14__out_11),
    .out_12(lb1d_14__out_12),
    .out_13(lb1d_14__out_13),
    .out_14(lb1d_14__out_14),
    .out_15(lb1d_14__out_15),
    .out_16(lb1d_14__out_16),
    .out_17(lb1d_14__out_17),
    .out_18(lb1d_14__out_18),
    .out_19(lb1d_14__out_19),
    .out_2(lb1d_14__out_2),
    .out_3(lb1d_14__out_3),
    .out_4(lb1d_14__out_4),
    .out_5(lb1d_14__out_5),
    .out_6(lb1d_14__out_6),
    .out_7(lb1d_14__out_7),
    .out_8(lb1d_14__out_8),
    .out_9(lb1d_14__out_9),
    .valid(lb1d_14__valid),
    .valid_chain(lb1d_14__valid_chain),
    .wen(lb1d_14__wen)
  );

  //Wire declarations for instance 'lb1d_15' (Module linebuffer_U3)
  wire  lb1d_15__clk;
  wire [15:0] lb1d_15__in_0;
  wire [15:0] lb1d_15__out_0;
  wire [15:0] lb1d_15__out_1;
  wire [15:0] lb1d_15__out_10;
  wire [15:0] lb1d_15__out_11;
  wire [15:0] lb1d_15__out_12;
  wire [15:0] lb1d_15__out_13;
  wire [15:0] lb1d_15__out_14;
  wire [15:0] lb1d_15__out_15;
  wire [15:0] lb1d_15__out_16;
  wire [15:0] lb1d_15__out_17;
  wire [15:0] lb1d_15__out_18;
  wire [15:0] lb1d_15__out_19;
  wire [15:0] lb1d_15__out_2;
  wire [15:0] lb1d_15__out_3;
  wire [15:0] lb1d_15__out_4;
  wire [15:0] lb1d_15__out_5;
  wire [15:0] lb1d_15__out_6;
  wire [15:0] lb1d_15__out_7;
  wire [15:0] lb1d_15__out_8;
  wire [15:0] lb1d_15__out_9;
  wire  lb1d_15__valid;
  wire  lb1d_15__valid_chain;
  wire  lb1d_15__wen;
  linebuffer_U3 lb1d_15(
    .clk(lb1d_15__clk),
    .in_0(lb1d_15__in_0),
    .out_0(lb1d_15__out_0),
    .out_1(lb1d_15__out_1),
    .out_10(lb1d_15__out_10),
    .out_11(lb1d_15__out_11),
    .out_12(lb1d_15__out_12),
    .out_13(lb1d_15__out_13),
    .out_14(lb1d_15__out_14),
    .out_15(lb1d_15__out_15),
    .out_16(lb1d_15__out_16),
    .out_17(lb1d_15__out_17),
    .out_18(lb1d_15__out_18),
    .out_19(lb1d_15__out_19),
    .out_2(lb1d_15__out_2),
    .out_3(lb1d_15__out_3),
    .out_4(lb1d_15__out_4),
    .out_5(lb1d_15__out_5),
    .out_6(lb1d_15__out_6),
    .out_7(lb1d_15__out_7),
    .out_8(lb1d_15__out_8),
    .out_9(lb1d_15__out_9),
    .valid(lb1d_15__valid),
    .valid_chain(lb1d_15__valid_chain),
    .wen(lb1d_15__wen)
  );

  //Wire declarations for instance 'lb1d_2' (Module linebuffer_U3)
  wire  lb1d_2__clk;
  wire [15:0] lb1d_2__in_0;
  wire [15:0] lb1d_2__out_0;
  wire [15:0] lb1d_2__out_1;
  wire [15:0] lb1d_2__out_10;
  wire [15:0] lb1d_2__out_11;
  wire [15:0] lb1d_2__out_12;
  wire [15:0] lb1d_2__out_13;
  wire [15:0] lb1d_2__out_14;
  wire [15:0] lb1d_2__out_15;
  wire [15:0] lb1d_2__out_16;
  wire [15:0] lb1d_2__out_17;
  wire [15:0] lb1d_2__out_18;
  wire [15:0] lb1d_2__out_19;
  wire [15:0] lb1d_2__out_2;
  wire [15:0] lb1d_2__out_3;
  wire [15:0] lb1d_2__out_4;
  wire [15:0] lb1d_2__out_5;
  wire [15:0] lb1d_2__out_6;
  wire [15:0] lb1d_2__out_7;
  wire [15:0] lb1d_2__out_8;
  wire [15:0] lb1d_2__out_9;
  wire  lb1d_2__valid;
  wire  lb1d_2__valid_chain;
  wire  lb1d_2__wen;
  linebuffer_U3 lb1d_2(
    .clk(lb1d_2__clk),
    .in_0(lb1d_2__in_0),
    .out_0(lb1d_2__out_0),
    .out_1(lb1d_2__out_1),
    .out_10(lb1d_2__out_10),
    .out_11(lb1d_2__out_11),
    .out_12(lb1d_2__out_12),
    .out_13(lb1d_2__out_13),
    .out_14(lb1d_2__out_14),
    .out_15(lb1d_2__out_15),
    .out_16(lb1d_2__out_16),
    .out_17(lb1d_2__out_17),
    .out_18(lb1d_2__out_18),
    .out_19(lb1d_2__out_19),
    .out_2(lb1d_2__out_2),
    .out_3(lb1d_2__out_3),
    .out_4(lb1d_2__out_4),
    .out_5(lb1d_2__out_5),
    .out_6(lb1d_2__out_6),
    .out_7(lb1d_2__out_7),
    .out_8(lb1d_2__out_8),
    .out_9(lb1d_2__out_9),
    .valid(lb1d_2__valid),
    .valid_chain(lb1d_2__valid_chain),
    .wen(lb1d_2__wen)
  );

  //Wire declarations for instance 'lb1d_3' (Module linebuffer_U3)
  wire  lb1d_3__clk;
  wire [15:0] lb1d_3__in_0;
  wire [15:0] lb1d_3__out_0;
  wire [15:0] lb1d_3__out_1;
  wire [15:0] lb1d_3__out_10;
  wire [15:0] lb1d_3__out_11;
  wire [15:0] lb1d_3__out_12;
  wire [15:0] lb1d_3__out_13;
  wire [15:0] lb1d_3__out_14;
  wire [15:0] lb1d_3__out_15;
  wire [15:0] lb1d_3__out_16;
  wire [15:0] lb1d_3__out_17;
  wire [15:0] lb1d_3__out_18;
  wire [15:0] lb1d_3__out_19;
  wire [15:0] lb1d_3__out_2;
  wire [15:0] lb1d_3__out_3;
  wire [15:0] lb1d_3__out_4;
  wire [15:0] lb1d_3__out_5;
  wire [15:0] lb1d_3__out_6;
  wire [15:0] lb1d_3__out_7;
  wire [15:0] lb1d_3__out_8;
  wire [15:0] lb1d_3__out_9;
  wire  lb1d_3__valid;
  wire  lb1d_3__valid_chain;
  wire  lb1d_3__wen;
  linebuffer_U3 lb1d_3(
    .clk(lb1d_3__clk),
    .in_0(lb1d_3__in_0),
    .out_0(lb1d_3__out_0),
    .out_1(lb1d_3__out_1),
    .out_10(lb1d_3__out_10),
    .out_11(lb1d_3__out_11),
    .out_12(lb1d_3__out_12),
    .out_13(lb1d_3__out_13),
    .out_14(lb1d_3__out_14),
    .out_15(lb1d_3__out_15),
    .out_16(lb1d_3__out_16),
    .out_17(lb1d_3__out_17),
    .out_18(lb1d_3__out_18),
    .out_19(lb1d_3__out_19),
    .out_2(lb1d_3__out_2),
    .out_3(lb1d_3__out_3),
    .out_4(lb1d_3__out_4),
    .out_5(lb1d_3__out_5),
    .out_6(lb1d_3__out_6),
    .out_7(lb1d_3__out_7),
    .out_8(lb1d_3__out_8),
    .out_9(lb1d_3__out_9),
    .valid(lb1d_3__valid),
    .valid_chain(lb1d_3__valid_chain),
    .wen(lb1d_3__wen)
  );

  //Wire declarations for instance 'lb1d_4' (Module linebuffer_U3)
  wire  lb1d_4__clk;
  wire [15:0] lb1d_4__in_0;
  wire [15:0] lb1d_4__out_0;
  wire [15:0] lb1d_4__out_1;
  wire [15:0] lb1d_4__out_10;
  wire [15:0] lb1d_4__out_11;
  wire [15:0] lb1d_4__out_12;
  wire [15:0] lb1d_4__out_13;
  wire [15:0] lb1d_4__out_14;
  wire [15:0] lb1d_4__out_15;
  wire [15:0] lb1d_4__out_16;
  wire [15:0] lb1d_4__out_17;
  wire [15:0] lb1d_4__out_18;
  wire [15:0] lb1d_4__out_19;
  wire [15:0] lb1d_4__out_2;
  wire [15:0] lb1d_4__out_3;
  wire [15:0] lb1d_4__out_4;
  wire [15:0] lb1d_4__out_5;
  wire [15:0] lb1d_4__out_6;
  wire [15:0] lb1d_4__out_7;
  wire [15:0] lb1d_4__out_8;
  wire [15:0] lb1d_4__out_9;
  wire  lb1d_4__valid;
  wire  lb1d_4__valid_chain;
  wire  lb1d_4__wen;
  linebuffer_U3 lb1d_4(
    .clk(lb1d_4__clk),
    .in_0(lb1d_4__in_0),
    .out_0(lb1d_4__out_0),
    .out_1(lb1d_4__out_1),
    .out_10(lb1d_4__out_10),
    .out_11(lb1d_4__out_11),
    .out_12(lb1d_4__out_12),
    .out_13(lb1d_4__out_13),
    .out_14(lb1d_4__out_14),
    .out_15(lb1d_4__out_15),
    .out_16(lb1d_4__out_16),
    .out_17(lb1d_4__out_17),
    .out_18(lb1d_4__out_18),
    .out_19(lb1d_4__out_19),
    .out_2(lb1d_4__out_2),
    .out_3(lb1d_4__out_3),
    .out_4(lb1d_4__out_4),
    .out_5(lb1d_4__out_5),
    .out_6(lb1d_4__out_6),
    .out_7(lb1d_4__out_7),
    .out_8(lb1d_4__out_8),
    .out_9(lb1d_4__out_9),
    .valid(lb1d_4__valid),
    .valid_chain(lb1d_4__valid_chain),
    .wen(lb1d_4__wen)
  );

  //Wire declarations for instance 'lb1d_5' (Module linebuffer_U3)
  wire  lb1d_5__clk;
  wire [15:0] lb1d_5__in_0;
  wire [15:0] lb1d_5__out_0;
  wire [15:0] lb1d_5__out_1;
  wire [15:0] lb1d_5__out_10;
  wire [15:0] lb1d_5__out_11;
  wire [15:0] lb1d_5__out_12;
  wire [15:0] lb1d_5__out_13;
  wire [15:0] lb1d_5__out_14;
  wire [15:0] lb1d_5__out_15;
  wire [15:0] lb1d_5__out_16;
  wire [15:0] lb1d_5__out_17;
  wire [15:0] lb1d_5__out_18;
  wire [15:0] lb1d_5__out_19;
  wire [15:0] lb1d_5__out_2;
  wire [15:0] lb1d_5__out_3;
  wire [15:0] lb1d_5__out_4;
  wire [15:0] lb1d_5__out_5;
  wire [15:0] lb1d_5__out_6;
  wire [15:0] lb1d_5__out_7;
  wire [15:0] lb1d_5__out_8;
  wire [15:0] lb1d_5__out_9;
  wire  lb1d_5__valid;
  wire  lb1d_5__valid_chain;
  wire  lb1d_5__wen;
  linebuffer_U3 lb1d_5(
    .clk(lb1d_5__clk),
    .in_0(lb1d_5__in_0),
    .out_0(lb1d_5__out_0),
    .out_1(lb1d_5__out_1),
    .out_10(lb1d_5__out_10),
    .out_11(lb1d_5__out_11),
    .out_12(lb1d_5__out_12),
    .out_13(lb1d_5__out_13),
    .out_14(lb1d_5__out_14),
    .out_15(lb1d_5__out_15),
    .out_16(lb1d_5__out_16),
    .out_17(lb1d_5__out_17),
    .out_18(lb1d_5__out_18),
    .out_19(lb1d_5__out_19),
    .out_2(lb1d_5__out_2),
    .out_3(lb1d_5__out_3),
    .out_4(lb1d_5__out_4),
    .out_5(lb1d_5__out_5),
    .out_6(lb1d_5__out_6),
    .out_7(lb1d_5__out_7),
    .out_8(lb1d_5__out_8),
    .out_9(lb1d_5__out_9),
    .valid(lb1d_5__valid),
    .valid_chain(lb1d_5__valid_chain),
    .wen(lb1d_5__wen)
  );

  //Wire declarations for instance 'lb1d_6' (Module linebuffer_U3)
  wire  lb1d_6__clk;
  wire [15:0] lb1d_6__in_0;
  wire [15:0] lb1d_6__out_0;
  wire [15:0] lb1d_6__out_1;
  wire [15:0] lb1d_6__out_10;
  wire [15:0] lb1d_6__out_11;
  wire [15:0] lb1d_6__out_12;
  wire [15:0] lb1d_6__out_13;
  wire [15:0] lb1d_6__out_14;
  wire [15:0] lb1d_6__out_15;
  wire [15:0] lb1d_6__out_16;
  wire [15:0] lb1d_6__out_17;
  wire [15:0] lb1d_6__out_18;
  wire [15:0] lb1d_6__out_19;
  wire [15:0] lb1d_6__out_2;
  wire [15:0] lb1d_6__out_3;
  wire [15:0] lb1d_6__out_4;
  wire [15:0] lb1d_6__out_5;
  wire [15:0] lb1d_6__out_6;
  wire [15:0] lb1d_6__out_7;
  wire [15:0] lb1d_6__out_8;
  wire [15:0] lb1d_6__out_9;
  wire  lb1d_6__valid;
  wire  lb1d_6__valid_chain;
  wire  lb1d_6__wen;
  linebuffer_U3 lb1d_6(
    .clk(lb1d_6__clk),
    .in_0(lb1d_6__in_0),
    .out_0(lb1d_6__out_0),
    .out_1(lb1d_6__out_1),
    .out_10(lb1d_6__out_10),
    .out_11(lb1d_6__out_11),
    .out_12(lb1d_6__out_12),
    .out_13(lb1d_6__out_13),
    .out_14(lb1d_6__out_14),
    .out_15(lb1d_6__out_15),
    .out_16(lb1d_6__out_16),
    .out_17(lb1d_6__out_17),
    .out_18(lb1d_6__out_18),
    .out_19(lb1d_6__out_19),
    .out_2(lb1d_6__out_2),
    .out_3(lb1d_6__out_3),
    .out_4(lb1d_6__out_4),
    .out_5(lb1d_6__out_5),
    .out_6(lb1d_6__out_6),
    .out_7(lb1d_6__out_7),
    .out_8(lb1d_6__out_8),
    .out_9(lb1d_6__out_9),
    .valid(lb1d_6__valid),
    .valid_chain(lb1d_6__valid_chain),
    .wen(lb1d_6__wen)
  );

  //Wire declarations for instance 'lb1d_7' (Module linebuffer_U3)
  wire  lb1d_7__clk;
  wire [15:0] lb1d_7__in_0;
  wire [15:0] lb1d_7__out_0;
  wire [15:0] lb1d_7__out_1;
  wire [15:0] lb1d_7__out_10;
  wire [15:0] lb1d_7__out_11;
  wire [15:0] lb1d_7__out_12;
  wire [15:0] lb1d_7__out_13;
  wire [15:0] lb1d_7__out_14;
  wire [15:0] lb1d_7__out_15;
  wire [15:0] lb1d_7__out_16;
  wire [15:0] lb1d_7__out_17;
  wire [15:0] lb1d_7__out_18;
  wire [15:0] lb1d_7__out_19;
  wire [15:0] lb1d_7__out_2;
  wire [15:0] lb1d_7__out_3;
  wire [15:0] lb1d_7__out_4;
  wire [15:0] lb1d_7__out_5;
  wire [15:0] lb1d_7__out_6;
  wire [15:0] lb1d_7__out_7;
  wire [15:0] lb1d_7__out_8;
  wire [15:0] lb1d_7__out_9;
  wire  lb1d_7__valid;
  wire  lb1d_7__valid_chain;
  wire  lb1d_7__wen;
  linebuffer_U3 lb1d_7(
    .clk(lb1d_7__clk),
    .in_0(lb1d_7__in_0),
    .out_0(lb1d_7__out_0),
    .out_1(lb1d_7__out_1),
    .out_10(lb1d_7__out_10),
    .out_11(lb1d_7__out_11),
    .out_12(lb1d_7__out_12),
    .out_13(lb1d_7__out_13),
    .out_14(lb1d_7__out_14),
    .out_15(lb1d_7__out_15),
    .out_16(lb1d_7__out_16),
    .out_17(lb1d_7__out_17),
    .out_18(lb1d_7__out_18),
    .out_19(lb1d_7__out_19),
    .out_2(lb1d_7__out_2),
    .out_3(lb1d_7__out_3),
    .out_4(lb1d_7__out_4),
    .out_5(lb1d_7__out_5),
    .out_6(lb1d_7__out_6),
    .out_7(lb1d_7__out_7),
    .out_8(lb1d_7__out_8),
    .out_9(lb1d_7__out_9),
    .valid(lb1d_7__valid),
    .valid_chain(lb1d_7__valid_chain),
    .wen(lb1d_7__wen)
  );

  //Wire declarations for instance 'lb1d_8' (Module linebuffer_U3)
  wire  lb1d_8__clk;
  wire [15:0] lb1d_8__in_0;
  wire [15:0] lb1d_8__out_0;
  wire [15:0] lb1d_8__out_1;
  wire [15:0] lb1d_8__out_10;
  wire [15:0] lb1d_8__out_11;
  wire [15:0] lb1d_8__out_12;
  wire [15:0] lb1d_8__out_13;
  wire [15:0] lb1d_8__out_14;
  wire [15:0] lb1d_8__out_15;
  wire [15:0] lb1d_8__out_16;
  wire [15:0] lb1d_8__out_17;
  wire [15:0] lb1d_8__out_18;
  wire [15:0] lb1d_8__out_19;
  wire [15:0] lb1d_8__out_2;
  wire [15:0] lb1d_8__out_3;
  wire [15:0] lb1d_8__out_4;
  wire [15:0] lb1d_8__out_5;
  wire [15:0] lb1d_8__out_6;
  wire [15:0] lb1d_8__out_7;
  wire [15:0] lb1d_8__out_8;
  wire [15:0] lb1d_8__out_9;
  wire  lb1d_8__valid;
  wire  lb1d_8__valid_chain;
  wire  lb1d_8__wen;
  linebuffer_U3 lb1d_8(
    .clk(lb1d_8__clk),
    .in_0(lb1d_8__in_0),
    .out_0(lb1d_8__out_0),
    .out_1(lb1d_8__out_1),
    .out_10(lb1d_8__out_10),
    .out_11(lb1d_8__out_11),
    .out_12(lb1d_8__out_12),
    .out_13(lb1d_8__out_13),
    .out_14(lb1d_8__out_14),
    .out_15(lb1d_8__out_15),
    .out_16(lb1d_8__out_16),
    .out_17(lb1d_8__out_17),
    .out_18(lb1d_8__out_18),
    .out_19(lb1d_8__out_19),
    .out_2(lb1d_8__out_2),
    .out_3(lb1d_8__out_3),
    .out_4(lb1d_8__out_4),
    .out_5(lb1d_8__out_5),
    .out_6(lb1d_8__out_6),
    .out_7(lb1d_8__out_7),
    .out_8(lb1d_8__out_8),
    .out_9(lb1d_8__out_9),
    .valid(lb1d_8__valid),
    .valid_chain(lb1d_8__valid_chain),
    .wen(lb1d_8__wen)
  );

  //Wire declarations for instance 'lb1d_9' (Module linebuffer_U3)
  wire  lb1d_9__clk;
  wire [15:0] lb1d_9__in_0;
  wire [15:0] lb1d_9__out_0;
  wire [15:0] lb1d_9__out_1;
  wire [15:0] lb1d_9__out_10;
  wire [15:0] lb1d_9__out_11;
  wire [15:0] lb1d_9__out_12;
  wire [15:0] lb1d_9__out_13;
  wire [15:0] lb1d_9__out_14;
  wire [15:0] lb1d_9__out_15;
  wire [15:0] lb1d_9__out_16;
  wire [15:0] lb1d_9__out_17;
  wire [15:0] lb1d_9__out_18;
  wire [15:0] lb1d_9__out_19;
  wire [15:0] lb1d_9__out_2;
  wire [15:0] lb1d_9__out_3;
  wire [15:0] lb1d_9__out_4;
  wire [15:0] lb1d_9__out_5;
  wire [15:0] lb1d_9__out_6;
  wire [15:0] lb1d_9__out_7;
  wire [15:0] lb1d_9__out_8;
  wire [15:0] lb1d_9__out_9;
  wire  lb1d_9__valid;
  wire  lb1d_9__valid_chain;
  wire  lb1d_9__wen;
  linebuffer_U3 lb1d_9(
    .clk(lb1d_9__clk),
    .in_0(lb1d_9__in_0),
    .out_0(lb1d_9__out_0),
    .out_1(lb1d_9__out_1),
    .out_10(lb1d_9__out_10),
    .out_11(lb1d_9__out_11),
    .out_12(lb1d_9__out_12),
    .out_13(lb1d_9__out_13),
    .out_14(lb1d_9__out_14),
    .out_15(lb1d_9__out_15),
    .out_16(lb1d_9__out_16),
    .out_17(lb1d_9__out_17),
    .out_18(lb1d_9__out_18),
    .out_19(lb1d_9__out_19),
    .out_2(lb1d_9__out_2),
    .out_3(lb1d_9__out_3),
    .out_4(lb1d_9__out_4),
    .out_5(lb1d_9__out_5),
    .out_6(lb1d_9__out_6),
    .out_7(lb1d_9__out_7),
    .out_8(lb1d_9__out_8),
    .out_9(lb1d_9__out_9),
    .valid(lb1d_9__valid),
    .valid_chain(lb1d_9__valid_chain),
    .wen(lb1d_9__wen)
  );

  //Wire declarations for instance 'lbmem_10_0' (Module rowbuffer_U4)
  wire  lbmem_10_0__clk;
  wire  lbmem_10_0__flush;
  wire [15:0] lbmem_10_0__rdata;
  wire  lbmem_10_0__valid;
  wire [15:0] lbmem_10_0__wdata;
  wire  lbmem_10_0__wen;
  rowbuffer_U4 lbmem_10_0(
    .clk(lbmem_10_0__clk),
    .flush(lbmem_10_0__flush),
    .rdata(lbmem_10_0__rdata),
    .valid(lbmem_10_0__valid),
    .wdata(lbmem_10_0__wdata),
    .wen(lbmem_10_0__wen)
  );

  //Wire declarations for instance 'lbmem_10_0_flush' (Module corebit_const)
  wire  lbmem_10_0_flush__out;
  corebit_const #(.value(0)) lbmem_10_0_flush(
    .out(lbmem_10_0_flush__out)
  );

  //Wire declarations for instance 'lbmem_11_0' (Module rowbuffer_U4)
  wire  lbmem_11_0__clk;
  wire  lbmem_11_0__flush;
  wire [15:0] lbmem_11_0__rdata;
  wire  lbmem_11_0__valid;
  wire [15:0] lbmem_11_0__wdata;
  wire  lbmem_11_0__wen;
  rowbuffer_U4 lbmem_11_0(
    .clk(lbmem_11_0__clk),
    .flush(lbmem_11_0__flush),
    .rdata(lbmem_11_0__rdata),
    .valid(lbmem_11_0__valid),
    .wdata(lbmem_11_0__wdata),
    .wen(lbmem_11_0__wen)
  );

  //Wire declarations for instance 'lbmem_11_0_flush' (Module corebit_const)
  wire  lbmem_11_0_flush__out;
  corebit_const #(.value(0)) lbmem_11_0_flush(
    .out(lbmem_11_0_flush__out)
  );

  //Wire declarations for instance 'lbmem_12_0' (Module rowbuffer_U4)
  wire  lbmem_12_0__clk;
  wire  lbmem_12_0__flush;
  wire [15:0] lbmem_12_0__rdata;
  wire  lbmem_12_0__valid;
  wire [15:0] lbmem_12_0__wdata;
  wire  lbmem_12_0__wen;
  rowbuffer_U4 lbmem_12_0(
    .clk(lbmem_12_0__clk),
    .flush(lbmem_12_0__flush),
    .rdata(lbmem_12_0__rdata),
    .valid(lbmem_12_0__valid),
    .wdata(lbmem_12_0__wdata),
    .wen(lbmem_12_0__wen)
  );

  //Wire declarations for instance 'lbmem_12_0_flush' (Module corebit_const)
  wire  lbmem_12_0_flush__out;
  corebit_const #(.value(0)) lbmem_12_0_flush(
    .out(lbmem_12_0_flush__out)
  );

  //Wire declarations for instance 'lbmem_13_0' (Module rowbuffer_U4)
  wire  lbmem_13_0__clk;
  wire  lbmem_13_0__flush;
  wire [15:0] lbmem_13_0__rdata;
  wire  lbmem_13_0__valid;
  wire [15:0] lbmem_13_0__wdata;
  wire  lbmem_13_0__wen;
  rowbuffer_U4 lbmem_13_0(
    .clk(lbmem_13_0__clk),
    .flush(lbmem_13_0__flush),
    .rdata(lbmem_13_0__rdata),
    .valid(lbmem_13_0__valid),
    .wdata(lbmem_13_0__wdata),
    .wen(lbmem_13_0__wen)
  );

  //Wire declarations for instance 'lbmem_13_0_flush' (Module corebit_const)
  wire  lbmem_13_0_flush__out;
  corebit_const #(.value(0)) lbmem_13_0_flush(
    .out(lbmem_13_0_flush__out)
  );

  //Wire declarations for instance 'lbmem_14_0' (Module rowbuffer_U4)
  wire  lbmem_14_0__clk;
  wire  lbmem_14_0__flush;
  wire [15:0] lbmem_14_0__rdata;
  wire  lbmem_14_0__valid;
  wire [15:0] lbmem_14_0__wdata;
  wire  lbmem_14_0__wen;
  rowbuffer_U4 lbmem_14_0(
    .clk(lbmem_14_0__clk),
    .flush(lbmem_14_0__flush),
    .rdata(lbmem_14_0__rdata),
    .valid(lbmem_14_0__valid),
    .wdata(lbmem_14_0__wdata),
    .wen(lbmem_14_0__wen)
  );

  //Wire declarations for instance 'lbmem_14_0_flush' (Module corebit_const)
  wire  lbmem_14_0_flush__out;
  corebit_const #(.value(0)) lbmem_14_0_flush(
    .out(lbmem_14_0_flush__out)
  );

  //Wire declarations for instance 'lbmem_15_0' (Module rowbuffer_U4)
  wire  lbmem_15_0__clk;
  wire  lbmem_15_0__flush;
  wire [15:0] lbmem_15_0__rdata;
  wire  lbmem_15_0__valid;
  wire [15:0] lbmem_15_0__wdata;
  wire  lbmem_15_0__wen;
  rowbuffer_U4 lbmem_15_0(
    .clk(lbmem_15_0__clk),
    .flush(lbmem_15_0__flush),
    .rdata(lbmem_15_0__rdata),
    .valid(lbmem_15_0__valid),
    .wdata(lbmem_15_0__wdata),
    .wen(lbmem_15_0__wen)
  );

  //Wire declarations for instance 'lbmem_15_0_flush' (Module corebit_const)
  wire  lbmem_15_0_flush__out;
  corebit_const #(.value(0)) lbmem_15_0_flush(
    .out(lbmem_15_0_flush__out)
  );

  //Wire declarations for instance 'lbmem_1_0' (Module rowbuffer_U4)
  wire  lbmem_1_0__clk;
  wire  lbmem_1_0__flush;
  wire [15:0] lbmem_1_0__rdata;
  wire  lbmem_1_0__valid;
  wire [15:0] lbmem_1_0__wdata;
  wire  lbmem_1_0__wen;
  rowbuffer_U4 lbmem_1_0(
    .clk(lbmem_1_0__clk),
    .flush(lbmem_1_0__flush),
    .rdata(lbmem_1_0__rdata),
    .valid(lbmem_1_0__valid),
    .wdata(lbmem_1_0__wdata),
    .wen(lbmem_1_0__wen)
  );

  //Wire declarations for instance 'lbmem_1_0_flush' (Module corebit_const)
  wire  lbmem_1_0_flush__out;
  corebit_const #(.value(0)) lbmem_1_0_flush(
    .out(lbmem_1_0_flush__out)
  );

  //Wire declarations for instance 'lbmem_2_0' (Module rowbuffer_U4)
  wire  lbmem_2_0__clk;
  wire  lbmem_2_0__flush;
  wire [15:0] lbmem_2_0__rdata;
  wire  lbmem_2_0__valid;
  wire [15:0] lbmem_2_0__wdata;
  wire  lbmem_2_0__wen;
  rowbuffer_U4 lbmem_2_0(
    .clk(lbmem_2_0__clk),
    .flush(lbmem_2_0__flush),
    .rdata(lbmem_2_0__rdata),
    .valid(lbmem_2_0__valid),
    .wdata(lbmem_2_0__wdata),
    .wen(lbmem_2_0__wen)
  );

  //Wire declarations for instance 'lbmem_2_0_flush' (Module corebit_const)
  wire  lbmem_2_0_flush__out;
  corebit_const #(.value(0)) lbmem_2_0_flush(
    .out(lbmem_2_0_flush__out)
  );

  //Wire declarations for instance 'lbmem_3_0' (Module rowbuffer_U4)
  wire  lbmem_3_0__clk;
  wire  lbmem_3_0__flush;
  wire [15:0] lbmem_3_0__rdata;
  wire  lbmem_3_0__valid;
  wire [15:0] lbmem_3_0__wdata;
  wire  lbmem_3_0__wen;
  rowbuffer_U4 lbmem_3_0(
    .clk(lbmem_3_0__clk),
    .flush(lbmem_3_0__flush),
    .rdata(lbmem_3_0__rdata),
    .valid(lbmem_3_0__valid),
    .wdata(lbmem_3_0__wdata),
    .wen(lbmem_3_0__wen)
  );

  //Wire declarations for instance 'lbmem_3_0_flush' (Module corebit_const)
  wire  lbmem_3_0_flush__out;
  corebit_const #(.value(0)) lbmem_3_0_flush(
    .out(lbmem_3_0_flush__out)
  );

  //Wire declarations for instance 'lbmem_4_0' (Module rowbuffer_U4)
  wire  lbmem_4_0__clk;
  wire  lbmem_4_0__flush;
  wire [15:0] lbmem_4_0__rdata;
  wire  lbmem_4_0__valid;
  wire [15:0] lbmem_4_0__wdata;
  wire  lbmem_4_0__wen;
  rowbuffer_U4 lbmem_4_0(
    .clk(lbmem_4_0__clk),
    .flush(lbmem_4_0__flush),
    .rdata(lbmem_4_0__rdata),
    .valid(lbmem_4_0__valid),
    .wdata(lbmem_4_0__wdata),
    .wen(lbmem_4_0__wen)
  );

  //Wire declarations for instance 'lbmem_4_0_flush' (Module corebit_const)
  wire  lbmem_4_0_flush__out;
  corebit_const #(.value(0)) lbmem_4_0_flush(
    .out(lbmem_4_0_flush__out)
  );

  //Wire declarations for instance 'lbmem_5_0' (Module rowbuffer_U4)
  wire  lbmem_5_0__clk;
  wire  lbmem_5_0__flush;
  wire [15:0] lbmem_5_0__rdata;
  wire  lbmem_5_0__valid;
  wire [15:0] lbmem_5_0__wdata;
  wire  lbmem_5_0__wen;
  rowbuffer_U4 lbmem_5_0(
    .clk(lbmem_5_0__clk),
    .flush(lbmem_5_0__flush),
    .rdata(lbmem_5_0__rdata),
    .valid(lbmem_5_0__valid),
    .wdata(lbmem_5_0__wdata),
    .wen(lbmem_5_0__wen)
  );

  //Wire declarations for instance 'lbmem_5_0_flush' (Module corebit_const)
  wire  lbmem_5_0_flush__out;
  corebit_const #(.value(0)) lbmem_5_0_flush(
    .out(lbmem_5_0_flush__out)
  );

  //Wire declarations for instance 'lbmem_6_0' (Module rowbuffer_U4)
  wire  lbmem_6_0__clk;
  wire  lbmem_6_0__flush;
  wire [15:0] lbmem_6_0__rdata;
  wire  lbmem_6_0__valid;
  wire [15:0] lbmem_6_0__wdata;
  wire  lbmem_6_0__wen;
  rowbuffer_U4 lbmem_6_0(
    .clk(lbmem_6_0__clk),
    .flush(lbmem_6_0__flush),
    .rdata(lbmem_6_0__rdata),
    .valid(lbmem_6_0__valid),
    .wdata(lbmem_6_0__wdata),
    .wen(lbmem_6_0__wen)
  );

  //Wire declarations for instance 'lbmem_6_0_flush' (Module corebit_const)
  wire  lbmem_6_0_flush__out;
  corebit_const #(.value(0)) lbmem_6_0_flush(
    .out(lbmem_6_0_flush__out)
  );

  //Wire declarations for instance 'lbmem_7_0' (Module rowbuffer_U4)
  wire  lbmem_7_0__clk;
  wire  lbmem_7_0__flush;
  wire [15:0] lbmem_7_0__rdata;
  wire  lbmem_7_0__valid;
  wire [15:0] lbmem_7_0__wdata;
  wire  lbmem_7_0__wen;
  rowbuffer_U4 lbmem_7_0(
    .clk(lbmem_7_0__clk),
    .flush(lbmem_7_0__flush),
    .rdata(lbmem_7_0__rdata),
    .valid(lbmem_7_0__valid),
    .wdata(lbmem_7_0__wdata),
    .wen(lbmem_7_0__wen)
  );

  //Wire declarations for instance 'lbmem_7_0_flush' (Module corebit_const)
  wire  lbmem_7_0_flush__out;
  corebit_const #(.value(0)) lbmem_7_0_flush(
    .out(lbmem_7_0_flush__out)
  );

  //Wire declarations for instance 'lbmem_8_0' (Module rowbuffer_U4)
  wire  lbmem_8_0__clk;
  wire  lbmem_8_0__flush;
  wire [15:0] lbmem_8_0__rdata;
  wire  lbmem_8_0__valid;
  wire [15:0] lbmem_8_0__wdata;
  wire  lbmem_8_0__wen;
  rowbuffer_U4 lbmem_8_0(
    .clk(lbmem_8_0__clk),
    .flush(lbmem_8_0__flush),
    .rdata(lbmem_8_0__rdata),
    .valid(lbmem_8_0__valid),
    .wdata(lbmem_8_0__wdata),
    .wen(lbmem_8_0__wen)
  );

  //Wire declarations for instance 'lbmem_8_0_flush' (Module corebit_const)
  wire  lbmem_8_0_flush__out;
  corebit_const #(.value(0)) lbmem_8_0_flush(
    .out(lbmem_8_0_flush__out)
  );

  //Wire declarations for instance 'lbmem_9_0' (Module rowbuffer_U4)
  wire  lbmem_9_0__clk;
  wire  lbmem_9_0__flush;
  wire [15:0] lbmem_9_0__rdata;
  wire  lbmem_9_0__valid;
  wire [15:0] lbmem_9_0__wdata;
  wire  lbmem_9_0__wen;
  rowbuffer_U4 lbmem_9_0(
    .clk(lbmem_9_0__clk),
    .flush(lbmem_9_0__flush),
    .rdata(lbmem_9_0__rdata),
    .valid(lbmem_9_0__valid),
    .wdata(lbmem_9_0__wdata),
    .wen(lbmem_9_0__wen)
  );

  //Wire declarations for instance 'lbmem_9_0_flush' (Module corebit_const)
  wire  lbmem_9_0_flush__out;
  corebit_const #(.value(0)) lbmem_9_0_flush(
    .out(lbmem_9_0_flush__out)
  );

  //Wire declarations for instance 'valcompare_0' (Module coreir_ule)
  wire [15:0] valcompare_0__in0;
  wire [15:0] valcompare_0__in1;
  wire  valcompare_0__out;
  coreir_ule #(.width(16)) valcompare_0(
    .in0(valcompare_0__in0),
    .in1(valcompare_0__in1),
    .out(valcompare_0__out)
  );

  //Wire declarations for instance 'valcompare_1' (Module coreir_ule)
  wire [15:0] valcompare_1__in0;
  wire [15:0] valcompare_1__in1;
  wire  valcompare_1__out;
  coreir_ule #(.width(16)) valcompare_1(
    .in0(valcompare_1__in0),
    .in1(valcompare_1__in1),
    .out(valcompare_1__out)
  );

  //Wire declarations for instance 'valcounter_0' (Module counter_U7)
  wire  valcounter_0__clk;
  wire  valcounter_0__en;
  wire [15:0] valcounter_0__out;
  wire  valcounter_0__overflow;
  wire  valcounter_0__reset;
  counter_U7 valcounter_0(
    .clk(valcounter_0__clk),
    .en(valcounter_0__en),
    .out(valcounter_0__out),
    .overflow(valcounter_0__overflow),
    .reset(valcounter_0__reset)
  );

  //Wire declarations for instance 'valcounter_0_reset' (Module corebit_const)
  wire  valcounter_0_reset__out;
  corebit_const #(.value(0)) valcounter_0_reset(
    .out(valcounter_0_reset__out)
  );

  //Wire declarations for instance 'valcounter_1' (Module counter_U8)
  wire  valcounter_1__clk;
  wire  valcounter_1__en;
  wire [15:0] valcounter_1__out;
  wire  valcounter_1__overflow;
  wire  valcounter_1__reset;
  counter_U8 valcounter_1(
    .clk(valcounter_1__clk),
    .en(valcounter_1__en),
    .out(valcounter_1__out),
    .overflow(valcounter_1__overflow),
    .reset(valcounter_1__reset)
  );

  //Wire declarations for instance 'valcounter_1_reset' (Module corebit_const)
  wire  valcounter_1_reset__out;
  corebit_const #(.value(0)) valcounter_1_reset(
    .out(valcounter_1_reset__out)
  );

  //Wire declarations for instance 'valid_andr' (Module bitopn_U9)
  wire [2:0] valid_andr__in;
  wire  valid_andr__out;
  bitopn_U9 valid_andr(
    .in(valid_andr__in),
    .out(valid_andr__out)
  );

  //All the connections
  assign lbmem_1_0__wen = wen;
  assign lbmem_1_0__wdata[15:0] = in_0_0[15:0];
  assign lbmem_1_0__flush = lbmem_1_0_flush__out;
  assign valcounter_0__en = wen;
  assign valid_andr__in[0] = wen;
  assign lb1d_0__wen = wen;
  assign lb1d_3__wen = wen;
  assign lb1d_1__wen = wen;
  assign lb1d_2__wen = wen;
  assign lb1d_4__wen = wen;
  assign lb1d_5__wen = wen;
  assign lb1d_6__wen = wen;
  assign lb1d_7__wen = wen;
  assign lb1d_8__wen = wen;
  assign lb1d_9__wen = wen;
  assign lb1d_10__wen = wen;
  assign lb1d_11__wen = wen;
  assign lb1d_12__wen = wen;
  assign lb1d_13__wen = wen;
  assign lb1d_14__wen = wen;
  assign lb1d_15__wen = wen;
  assign lbmem_2_0__wdata[15:0] = lbmem_1_0__rdata[15:0];
  assign lb1d_1__in_0[15:0] = lbmem_1_0__rdata[15:0];
  assign lbmem_2_0__wen = lbmem_1_0__valid;
  assign lbmem_2_0__flush = lbmem_2_0_flush__out;
  assign lbmem_3_0__wdata[15:0] = lbmem_2_0__rdata[15:0];
  assign lb1d_2__in_0[15:0] = lbmem_2_0__rdata[15:0];
  assign lbmem_3_0__wen = lbmem_2_0__valid;
  assign lbmem_3_0__flush = lbmem_3_0_flush__out;
  assign lbmem_4_0__wdata[15:0] = lbmem_3_0__rdata[15:0];
  assign lb1d_3__in_0[15:0] = lbmem_3_0__rdata[15:0];
  assign lbmem_4_0__wen = lbmem_3_0__valid;
  assign lbmem_4_0__flush = lbmem_4_0_flush__out;
  assign lbmem_5_0__wdata[15:0] = lbmem_4_0__rdata[15:0];
  assign lb1d_4__in_0[15:0] = lbmem_4_0__rdata[15:0];
  assign lbmem_5_0__wen = lbmem_4_0__valid;
  assign lbmem_5_0__flush = lbmem_5_0_flush__out;
  assign lbmem_6_0__wdata[15:0] = lbmem_5_0__rdata[15:0];
  assign lb1d_5__in_0[15:0] = lbmem_5_0__rdata[15:0];
  assign lbmem_6_0__wen = lbmem_5_0__valid;
  assign lbmem_6_0__flush = lbmem_6_0_flush__out;
  assign lbmem_7_0__wdata[15:0] = lbmem_6_0__rdata[15:0];
  assign lb1d_6__in_0[15:0] = lbmem_6_0__rdata[15:0];
  assign lbmem_7_0__wen = lbmem_6_0__valid;
  assign lbmem_7_0__flush = lbmem_7_0_flush__out;
  assign lbmem_8_0__wdata[15:0] = lbmem_7_0__rdata[15:0];
  assign lb1d_7__in_0[15:0] = lbmem_7_0__rdata[15:0];
  assign lbmem_8_0__wen = lbmem_7_0__valid;
  assign lbmem_8_0__flush = lbmem_8_0_flush__out;
  assign lbmem_9_0__wdata[15:0] = lbmem_8_0__rdata[15:0];
  assign lb1d_8__in_0[15:0] = lbmem_8_0__rdata[15:0];
  assign lbmem_9_0__wen = lbmem_8_0__valid;
  assign lbmem_9_0__flush = lbmem_9_0_flush__out;
  assign lbmem_10_0__wdata[15:0] = lbmem_9_0__rdata[15:0];
  assign lb1d_9__in_0[15:0] = lbmem_9_0__rdata[15:0];
  assign lbmem_10_0__flush = lbmem_10_0_flush__out;
  assign lbmem_10_0__wen = lbmem_9_0__valid;
  assign lbmem_11_0__wdata[15:0] = lbmem_10_0__rdata[15:0];
  assign lb1d_10__in_0[15:0] = lbmem_10_0__rdata[15:0];
  assign lbmem_11_0__flush = lbmem_11_0_flush__out;
  assign lbmem_11_0__wen = lbmem_10_0__valid;
  assign lbmem_12_0__wdata[15:0] = lbmem_11_0__rdata[15:0];
  assign lb1d_11__in_0[15:0] = lbmem_11_0__rdata[15:0];
  assign lbmem_12_0__flush = lbmem_12_0_flush__out;
  assign lbmem_12_0__wen = lbmem_11_0__valid;
  assign lbmem_13_0__wdata[15:0] = lbmem_12_0__rdata[15:0];
  assign lb1d_12__in_0[15:0] = lbmem_12_0__rdata[15:0];
  assign lbmem_13_0__flush = lbmem_13_0_flush__out;
  assign lbmem_13_0__wen = lbmem_12_0__valid;
  assign lbmem_14_0__wdata[15:0] = lbmem_13_0__rdata[15:0];
  assign lb1d_13__in_0[15:0] = lbmem_13_0__rdata[15:0];
  assign lbmem_14_0__flush = lbmem_14_0_flush__out;
  assign lbmem_14_0__wen = lbmem_13_0__valid;
  assign lbmem_15_0__wdata[15:0] = lbmem_14_0__rdata[15:0];
  assign lb1d_14__in_0[15:0] = lbmem_14_0__rdata[15:0];
  assign lbmem_15_0__flush = lbmem_15_0_flush__out;
  assign lbmem_15_0__wen = lbmem_14_0__valid;
  assign lb1d_15__in_0[15:0] = lbmem_15_0__rdata[15:0];
  assign valid_chain = lbmem_15_0__valid;
  assign valcounter_0__reset = valcounter_0_reset__out;
  assign valcompare_0__in1[15:0] = valcounter_0__out[15:0];
  assign valcompare_0__in0[15:0] = const_stencil0__out[15:0];
  assign valcompare_1__in0[15:0] = const_stencil1__out[15:0];
  assign valcounter_1__reset = valcounter_1_reset__out;
  assign valcounter_1__en = valcounter_0__overflow;
  assign valcompare_1__in1[15:0] = valcounter_1__out[15:0];
  assign valid_andr__in[1] = valcompare_0__out;
  assign valid = valid_andr__out;
  assign valid_andr__in[2] = valcompare_1__out;
  assign out_15_0[15:0] = lb1d_0__out_0[15:0];
  assign out_1_7[15:0] = lb1d_14__out_7[15:0];
  assign out_15_10[15:0] = lb1d_0__out_10[15:0];
  assign out_2_4[15:0] = lb1d_13__out_4[15:0];
  assign lb1d_0__clk = clk;
  assign lb1d_1__clk = clk;
  assign lb1d_10__clk = clk;
  assign lb1d_11__clk = clk;
  assign lb1d_12__clk = clk;
  assign lb1d_13__clk = clk;
  assign lb1d_14__clk = clk;
  assign lb1d_15__clk = clk;
  assign lb1d_2__clk = clk;
  assign lb1d_3__clk = clk;
  assign lb1d_4__clk = clk;
  assign lb1d_5__clk = clk;
  assign lb1d_6__clk = clk;
  assign lb1d_7__clk = clk;
  assign lb1d_8__clk = clk;
  assign lb1d_9__clk = clk;
  assign lbmem_10_0__clk = clk;
  assign lbmem_11_0__clk = clk;
  assign lbmem_12_0__clk = clk;
  assign lbmem_13_0__clk = clk;
  assign lbmem_14_0__clk = clk;
  assign lbmem_15_0__clk = clk;
  assign lbmem_1_0__clk = clk;
  assign lbmem_2_0__clk = clk;
  assign lbmem_3_0__clk = clk;
  assign lbmem_4_0__clk = clk;
  assign lbmem_5_0__clk = clk;
  assign lbmem_6_0__clk = clk;
  assign lbmem_7_0__clk = clk;
  assign lbmem_8_0__clk = clk;
  assign lbmem_9_0__clk = clk;
  assign valcounter_0__clk = clk;
  assign valcounter_1__clk = clk;
  assign out_4_4[15:0] = lb1d_11__out_4[15:0];
  assign out_13_5[15:0] = lb1d_2__out_5[15:0];
  assign out_4_12[15:0] = lb1d_11__out_12[15:0];
  assign out_15_12[15:0] = lb1d_0__out_12[15:0];
  assign out_4_2[15:0] = lb1d_11__out_2[15:0];
  assign out_15_1[15:0] = lb1d_0__out_1[15:0];
  assign out_5_4[15:0] = lb1d_10__out_4[15:0];
  assign out_15_2[15:0] = lb1d_0__out_2[15:0];
  assign out_0_7[15:0] = lb1d_15__out_7[15:0];
  assign out_15_3[15:0] = lb1d_0__out_3[15:0];
  assign out_15_4[15:0] = lb1d_0__out_4[15:0];
  assign out_11_1[15:0] = lb1d_4__out_1[15:0];
  assign out_15_5[15:0] = lb1d_0__out_5[15:0];
  assign out_7_0[15:0] = lb1d_8__out_0[15:0];
  assign out_15_6[15:0] = lb1d_0__out_6[15:0];
  assign out_5_0[15:0] = lb1d_10__out_0[15:0];
  assign out_15_7[15:0] = lb1d_0__out_7[15:0];
  assign out_3_0[15:0] = lb1d_12__out_0[15:0];
  assign out_15_8[15:0] = lb1d_0__out_8[15:0];
  assign out_0_2[15:0] = lb1d_15__out_2[15:0];
  assign out_15_9[15:0] = lb1d_0__out_9[15:0];
  assign out_5_1[15:0] = lb1d_10__out_1[15:0];
  assign out_4_3[15:0] = lb1d_11__out_3[15:0];
  assign out_15_11[15:0] = lb1d_0__out_11[15:0];
  assign out_10_6[15:0] = lb1d_5__out_6[15:0];
  assign lb1d_0__in_0[15:0] = in_0_0[15:0];
  assign out_4_1[15:0] = lb1d_11__out_1[15:0];
  assign out_2_8[15:0] = lb1d_13__out_8[15:0];
  assign out_14_7[15:0] = lb1d_1__out_7[15:0];
  assign out_1_6[15:0] = lb1d_14__out_6[15:0];
  assign out_14_8[15:0] = lb1d_1__out_8[15:0];
  assign out_5_6[15:0] = lb1d_10__out_6[15:0];
  assign out_3_6[15:0] = lb1d_12__out_6[15:0];
  assign out_14_3[15:0] = lb1d_1__out_3[15:0];
  assign out_2_3[15:0] = lb1d_13__out_3[15:0];
  assign out_14_4[15:0] = lb1d_1__out_4[15:0];
  assign out_14_5[15:0] = lb1d_1__out_5[15:0];
  assign out_13_0[15:0] = lb1d_2__out_0[15:0];
  assign out_14_6[15:0] = lb1d_1__out_6[15:0];
  assign out_0_4[15:0] = lb1d_15__out_4[15:0];
  assign out_3_2[15:0] = lb1d_12__out_2[15:0];
  assign out_4_7[15:0] = lb1d_11__out_7[15:0];
  assign out_14_0[15:0] = lb1d_1__out_0[15:0];
  assign out_1_8[15:0] = lb1d_14__out_8[15:0];
  assign out_3_3[15:0] = lb1d_12__out_3[15:0];
  assign out_14_1[15:0] = lb1d_1__out_1[15:0];
  assign out_1_1[15:0] = lb1d_14__out_1[15:0];
  assign out_14_2[15:0] = lb1d_1__out_2[15:0];
  assign out_3_5[15:0] = lb1d_12__out_5[15:0];
  assign out_14_9[15:0] = lb1d_1__out_9[15:0];
  assign out_4_0[15:0] = lb1d_11__out_0[15:0];
  assign out_13_4[15:0] = lb1d_2__out_4[15:0];
  assign out_5_3[15:0] = lb1d_10__out_3[15:0];
  assign out_5_5[15:0] = lb1d_10__out_5[15:0];
  assign out_4_8[15:0] = lb1d_11__out_8[15:0];
  assign out_15_13[15:0] = lb1d_0__out_13[15:0];
  assign out_4_6[15:0] = lb1d_11__out_6[15:0];
  assign out_15_14[15:0] = lb1d_0__out_14[15:0];
  assign out_14_11[15:0] = lb1d_1__out_11[15:0];
  assign out_15_15[15:0] = lb1d_0__out_15[15:0];
  assign out_7_1[15:0] = lb1d_8__out_1[15:0];
  assign out_15_16[15:0] = lb1d_0__out_16[15:0];
  assign out_15_17[15:0] = lb1d_0__out_17[15:0];
  assign out_4_5[15:0] = lb1d_11__out_5[15:0];
  assign out_15_18[15:0] = lb1d_0__out_18[15:0];
  assign out_2_0[15:0] = lb1d_13__out_0[15:0];
  assign out_15_19[15:0] = lb1d_0__out_19[15:0];
  assign out_11_3[15:0] = lb1d_4__out_3[15:0];
  assign out_14_12[15:0] = lb1d_1__out_12[15:0];
  assign out_5_2[15:0] = lb1d_10__out_2[15:0];
  assign out_2_7[15:0] = lb1d_13__out_7[15:0];
  assign out_3_4[15:0] = lb1d_12__out_4[15:0];
  assign out_14_10[15:0] = lb1d_1__out_10[15:0];
  assign out_14_13[15:0] = lb1d_1__out_13[15:0];
  assign out_14_14[15:0] = lb1d_1__out_14[15:0];
  assign out_5_8[15:0] = lb1d_10__out_8[15:0];
  assign out_14_15[15:0] = lb1d_1__out_15[15:0];
  assign out_9_2[15:0] = lb1d_6__out_2[15:0];
  assign out_14_16[15:0] = lb1d_1__out_16[15:0];
  assign out_5_9[15:0] = lb1d_10__out_9[15:0];
  assign out_14_17[15:0] = lb1d_1__out_17[15:0];
  assign out_14_18[15:0] = lb1d_1__out_18[15:0];
  assign out_5_10[15:0] = lb1d_10__out_10[15:0];
  assign out_14_19[15:0] = lb1d_1__out_19[15:0];
  assign out_2_5[15:0] = lb1d_13__out_5[15:0];
  assign out_1_2[15:0] = lb1d_14__out_2[15:0];
  assign out_5_11[15:0] = lb1d_10__out_11[15:0];
  assign out_5_7[15:0] = lb1d_10__out_7[15:0];
  assign out_5_12[15:0] = lb1d_10__out_12[15:0];
  assign out_4_9[15:0] = lb1d_11__out_9[15:0];
  assign out_5_13[15:0] = lb1d_10__out_13[15:0];
  assign out_2_1[15:0] = lb1d_13__out_1[15:0];
  assign out_5_14[15:0] = lb1d_10__out_14[15:0];
  assign out_4_10[15:0] = lb1d_11__out_10[15:0];
  assign out_5_15[15:0] = lb1d_10__out_15[15:0];
  assign out_9_1[15:0] = lb1d_6__out_1[15:0];
  assign out_5_16[15:0] = lb1d_10__out_16[15:0];
  assign out_4_11[15:0] = lb1d_11__out_11[15:0];
  assign out_5_17[15:0] = lb1d_10__out_17[15:0];
  assign out_11_2[15:0] = lb1d_4__out_2[15:0];
  assign out_5_18[15:0] = lb1d_10__out_18[15:0];
  assign out_2_6[15:0] = lb1d_13__out_6[15:0];
  assign out_5_19[15:0] = lb1d_10__out_19[15:0];
  assign out_0_3[15:0] = lb1d_15__out_3[15:0];
  assign out_0_6[15:0] = lb1d_15__out_6[15:0];
  assign out_8_0[15:0] = lb1d_7__out_0[15:0];
  assign out_0_8[15:0] = lb1d_15__out_8[15:0];
  assign out_3_1[15:0] = lb1d_12__out_1[15:0];
  assign out_1_9[15:0] = lb1d_14__out_9[15:0];
  assign out_4_13[15:0] = lb1d_11__out_13[15:0];
  assign out_3_7[15:0] = lb1d_12__out_7[15:0];
  assign out_4_14[15:0] = lb1d_11__out_14[15:0];
  assign out_1_3[15:0] = lb1d_14__out_3[15:0];
  assign out_4_15[15:0] = lb1d_11__out_15[15:0];
  assign out_3_8[15:0] = lb1d_12__out_8[15:0];
  assign out_4_16[15:0] = lb1d_11__out_16[15:0];
  assign out_4_17[15:0] = lb1d_11__out_17[15:0];
  assign out_3_9[15:0] = lb1d_12__out_9[15:0];
  assign out_4_18[15:0] = lb1d_11__out_18[15:0];
  assign out_1_4[15:0] = lb1d_14__out_4[15:0];
  assign out_4_19[15:0] = lb1d_11__out_19[15:0];
  assign out_3_11[15:0] = lb1d_12__out_11[15:0];
  assign out_3_10[15:0] = lb1d_12__out_10[15:0];
  assign out_2_2[15:0] = lb1d_13__out_2[15:0];
  assign out_0_1[15:0] = lb1d_15__out_1[15:0];
  assign out_2_9[15:0] = lb1d_13__out_9[15:0];
  assign out_3_12[15:0] = lb1d_12__out_12[15:0];
  assign out_0_9[15:0] = lb1d_15__out_9[15:0];
  assign out_3_13[15:0] = lb1d_12__out_13[15:0];
  assign out_13_3[15:0] = lb1d_2__out_3[15:0];
  assign out_3_14[15:0] = lb1d_12__out_14[15:0];
  assign out_3_15[15:0] = lb1d_12__out_15[15:0];
  assign out_12_1[15:0] = lb1d_3__out_1[15:0];
  assign out_3_16[15:0] = lb1d_12__out_16[15:0];
  assign out_10_7[15:0] = lb1d_5__out_7[15:0];
  assign out_3_17[15:0] = lb1d_12__out_17[15:0];
  assign out_1_0[15:0] = lb1d_14__out_0[15:0];
  assign out_3_18[15:0] = lb1d_12__out_18[15:0];
  assign out_13_1[15:0] = lb1d_2__out_1[15:0];
  assign out_3_19[15:0] = lb1d_12__out_19[15:0];
  assign out_12_2[15:0] = lb1d_3__out_2[15:0];
  assign out_2_10[15:0] = lb1d_13__out_10[15:0];
  assign out_1_5[15:0] = lb1d_14__out_5[15:0];
  assign out_11_5[15:0] = lb1d_4__out_5[15:0];
  assign out_2_11[15:0] = lb1d_13__out_11[15:0];
  assign out_13_2[15:0] = lb1d_2__out_2[15:0];
  assign out_0_11[15:0] = lb1d_15__out_11[15:0];
  assign out_2_12[15:0] = lb1d_13__out_12[15:0];
  assign out_10_3[15:0] = lb1d_5__out_3[15:0];
  assign out_2_13[15:0] = lb1d_13__out_13[15:0];
  assign out_8_4[15:0] = lb1d_7__out_4[15:0];
  assign out_2_14[15:0] = lb1d_13__out_14[15:0];
  assign out_2_15[15:0] = lb1d_13__out_15[15:0];
  assign out_2_16[15:0] = lb1d_13__out_16[15:0];
  assign out_12_6[15:0] = lb1d_3__out_6[15:0];
  assign out_2_17[15:0] = lb1d_13__out_17[15:0];
  assign out_0_0[15:0] = lb1d_15__out_0[15:0];
  assign out_2_18[15:0] = lb1d_13__out_18[15:0];
  assign out_10_9[15:0] = lb1d_5__out_9[15:0];
  assign out_2_19[15:0] = lb1d_13__out_19[15:0];
  assign out_8_5[15:0] = lb1d_7__out_5[15:0];
  assign out_1_10[15:0] = lb1d_14__out_10[15:0];
  assign out_0_5[15:0] = lb1d_15__out_5[15:0];
  assign out_7_5[15:0] = lb1d_8__out_5[15:0];
  assign out_1_11[15:0] = lb1d_14__out_11[15:0];
  assign out_1_12[15:0] = lb1d_14__out_12[15:0];
  assign out_0_10[15:0] = lb1d_15__out_10[15:0];
  assign out_1_13[15:0] = lb1d_14__out_13[15:0];
  assign out_8_1[15:0] = lb1d_7__out_1[15:0];
  assign out_1_14[15:0] = lb1d_14__out_14[15:0];
  assign out_1_15[15:0] = lb1d_14__out_15[15:0];
  assign out_12_3[15:0] = lb1d_3__out_3[15:0];
  assign out_1_16[15:0] = lb1d_14__out_16[15:0];
  assign out_1_17[15:0] = lb1d_14__out_17[15:0];
  assign out_12_4[15:0] = lb1d_3__out_4[15:0];
  assign out_1_18[15:0] = lb1d_14__out_18[15:0];
  assign out_8_7[15:0] = lb1d_7__out_7[15:0];
  assign out_1_19[15:0] = lb1d_14__out_19[15:0];
  assign out_10_0[15:0] = lb1d_5__out_0[15:0];
  assign out_12_5[15:0] = lb1d_3__out_5[15:0];
  assign out_13_6[15:0] = lb1d_2__out_6[15:0];
  assign out_11_6[15:0] = lb1d_4__out_6[15:0];
  assign out_10_4[15:0] = lb1d_5__out_4[15:0];
  assign out_13_7[15:0] = lb1d_2__out_7[15:0];
  assign out_0_12[15:0] = lb1d_15__out_12[15:0];
  assign out_0_13[15:0] = lb1d_15__out_13[15:0];
  assign out_13_8[15:0] = lb1d_2__out_8[15:0];
  assign out_0_14[15:0] = lb1d_15__out_14[15:0];
  assign out_8_2[15:0] = lb1d_7__out_2[15:0];
  assign out_0_15[15:0] = lb1d_15__out_15[15:0];
  assign out_13_9[15:0] = lb1d_2__out_9[15:0];
  assign out_0_16[15:0] = lb1d_15__out_16[15:0];
  assign out_9_6[15:0] = lb1d_6__out_6[15:0];
  assign out_0_17[15:0] = lb1d_15__out_17[15:0];
  assign out_13_10[15:0] = lb1d_2__out_10[15:0];
  assign out_0_18[15:0] = lb1d_15__out_18[15:0];
  assign out_11_4[15:0] = lb1d_4__out_4[15:0];
  assign out_0_19[15:0] = lb1d_15__out_19[15:0];
  assign out_10_5[15:0] = lb1d_5__out_5[15:0];
  assign out_13_11[15:0] = lb1d_2__out_11[15:0];
  assign out_12_0[15:0] = lb1d_3__out_0[15:0];
  assign out_7_3[15:0] = lb1d_8__out_3[15:0];
  assign out_12_7[15:0] = lb1d_3__out_7[15:0];
  assign out_6_6[15:0] = lb1d_9__out_6[15:0];
  assign out_13_12[15:0] = lb1d_2__out_12[15:0];
  assign out_13_13[15:0] = lb1d_2__out_13[15:0];
  assign out_12_8[15:0] = lb1d_3__out_8[15:0];
  assign out_13_14[15:0] = lb1d_2__out_14[15:0];
  assign out_13_15[15:0] = lb1d_2__out_15[15:0];
  assign out_12_9[15:0] = lb1d_3__out_9[15:0];
  assign out_13_16[15:0] = lb1d_2__out_16[15:0];
  assign out_10_1[15:0] = lb1d_5__out_1[15:0];
  assign out_13_17[15:0] = lb1d_2__out_17[15:0];
  assign out_12_10[15:0] = lb1d_3__out_10[15:0];
  assign out_13_18[15:0] = lb1d_2__out_18[15:0];
  assign out_10_8[15:0] = lb1d_5__out_8[15:0];
  assign out_13_19[15:0] = lb1d_2__out_19[15:0];
  assign out_12_11[15:0] = lb1d_3__out_11[15:0];
  assign out_9_8[15:0] = lb1d_6__out_8[15:0];
  assign out_11_0[15:0] = lb1d_4__out_0[15:0];
  assign out_12_12[15:0] = lb1d_3__out_12[15:0];
  assign out_12_13[15:0] = lb1d_3__out_13[15:0];
  assign out_11_7[15:0] = lb1d_4__out_7[15:0];
  assign out_12_14[15:0] = lb1d_3__out_14[15:0];
  assign out_9_3[15:0] = lb1d_6__out_3[15:0];
  assign out_12_15[15:0] = lb1d_3__out_15[15:0];
  assign out_11_8[15:0] = lb1d_4__out_8[15:0];
  assign out_12_16[15:0] = lb1d_3__out_16[15:0];
  assign out_12_17[15:0] = lb1d_3__out_17[15:0];
  assign out_11_9[15:0] = lb1d_4__out_9[15:0];
  assign out_12_18[15:0] = lb1d_3__out_18[15:0];
  assign out_9_4[15:0] = lb1d_6__out_4[15:0];
  assign out_12_19[15:0] = lb1d_3__out_19[15:0];
  assign out_11_10[15:0] = lb1d_4__out_10[15:0];
  assign out_9_7[15:0] = lb1d_6__out_7[15:0];
  assign out_11_11[15:0] = lb1d_4__out_11[15:0];
  assign out_10_2[15:0] = lb1d_5__out_2[15:0];
  assign out_10_10[15:0] = lb1d_5__out_10[15:0];
  assign out_11_12[15:0] = lb1d_4__out_12[15:0];
  assign out_11_13[15:0] = lb1d_4__out_13[15:0];
  assign out_7_2[15:0] = lb1d_8__out_2[15:0];
  assign out_11_14[15:0] = lb1d_4__out_14[15:0];
  assign out_11_15[15:0] = lb1d_4__out_15[15:0];
  assign out_6_2[15:0] = lb1d_9__out_2[15:0];
  assign out_11_16[15:0] = lb1d_4__out_16[15:0];
  assign out_6_1[15:0] = lb1d_9__out_1[15:0];
  assign out_11_17[15:0] = lb1d_4__out_17[15:0];
  assign out_9_0[15:0] = lb1d_6__out_0[15:0];
  assign out_11_18[15:0] = lb1d_4__out_18[15:0];
  assign out_11_19[15:0] = lb1d_4__out_19[15:0];
  assign out_9_9[15:0] = lb1d_6__out_9[15:0];
  assign out_9_5[15:0] = lb1d_6__out_5[15:0];
  assign out_10_11[15:0] = lb1d_5__out_11[15:0];
  assign out_8_10[15:0] = lb1d_7__out_10[15:0];
  assign out_10_12[15:0] = lb1d_5__out_12[15:0];
  assign out_9_10[15:0] = lb1d_6__out_10[15:0];
  assign out_10_13[15:0] = lb1d_5__out_13[15:0];
  assign out_8_6[15:0] = lb1d_7__out_6[15:0];
  assign out_10_14[15:0] = lb1d_5__out_14[15:0];
  assign out_7_4[15:0] = lb1d_8__out_4[15:0];
  assign out_10_15[15:0] = lb1d_5__out_15[15:0];
  assign out_10_16[15:0] = lb1d_5__out_16[15:0];
  assign out_10_17[15:0] = lb1d_5__out_17[15:0];
  assign out_10_18[15:0] = lb1d_5__out_18[15:0];
  assign out_10_19[15:0] = lb1d_5__out_19[15:0];
  assign out_8_8[15:0] = lb1d_7__out_8[15:0];
  assign out_8_12[15:0] = lb1d_7__out_12[15:0];
  assign out_8_3[15:0] = lb1d_7__out_3[15:0];
  assign out_9_11[15:0] = lb1d_6__out_11[15:0];
  assign out_7_6[15:0] = lb1d_8__out_6[15:0];
  assign out_8_9[15:0] = lb1d_7__out_9[15:0];
  assign out_9_12[15:0] = lb1d_6__out_12[15:0];
  assign out_9_13[15:0] = lb1d_6__out_13[15:0];
  assign out_9_14[15:0] = lb1d_6__out_14[15:0];
  assign out_6_3[15:0] = lb1d_9__out_3[15:0];
  assign out_9_15[15:0] = lb1d_6__out_15[15:0];
  assign out_9_16[15:0] = lb1d_6__out_16[15:0];
  assign out_6_4[15:0] = lb1d_9__out_4[15:0];
  assign out_9_17[15:0] = lb1d_6__out_17[15:0];
  assign out_6_5[15:0] = lb1d_9__out_5[15:0];
  assign out_9_18[15:0] = lb1d_6__out_18[15:0];
  assign out_9_19[15:0] = lb1d_6__out_19[15:0];
  assign out_8_11[15:0] = lb1d_7__out_11[15:0];
  assign out_7_7[15:0] = lb1d_8__out_7[15:0];
  assign out_8_13[15:0] = lb1d_7__out_13[15:0];
  assign out_7_8[15:0] = lb1d_8__out_8[15:0];
  assign out_8_14[15:0] = lb1d_7__out_14[15:0];
  assign out_8_15[15:0] = lb1d_7__out_15[15:0];
  assign out_7_9[15:0] = lb1d_8__out_9[15:0];
  assign out_8_16[15:0] = lb1d_7__out_16[15:0];
  assign out_8_17[15:0] = lb1d_7__out_17[15:0];
  assign out_7_10[15:0] = lb1d_8__out_10[15:0];
  assign out_8_18[15:0] = lb1d_7__out_18[15:0];
  assign out_8_19[15:0] = lb1d_7__out_19[15:0];
  assign out_7_11[15:0] = lb1d_8__out_11[15:0];
  assign out_6_0[15:0] = lb1d_9__out_0[15:0];
  assign out_6_7[15:0] = lb1d_9__out_7[15:0];
  assign out_7_12[15:0] = lb1d_8__out_12[15:0];
  assign out_7_13[15:0] = lb1d_8__out_13[15:0];
  assign out_6_8[15:0] = lb1d_9__out_8[15:0];
  assign out_7_14[15:0] = lb1d_8__out_14[15:0];
  assign out_7_15[15:0] = lb1d_8__out_15[15:0];
  assign out_6_9[15:0] = lb1d_9__out_9[15:0];
  assign out_7_16[15:0] = lb1d_8__out_16[15:0];
  assign out_7_17[15:0] = lb1d_8__out_17[15:0];
  assign out_6_10[15:0] = lb1d_9__out_10[15:0];
  assign out_7_18[15:0] = lb1d_8__out_18[15:0];
  assign out_7_19[15:0] = lb1d_8__out_19[15:0];
  assign out_6_11[15:0] = lb1d_9__out_11[15:0];
  assign out_6_12[15:0] = lb1d_9__out_12[15:0];
  assign out_6_13[15:0] = lb1d_9__out_13[15:0];
  assign out_6_14[15:0] = lb1d_9__out_14[15:0];
  assign out_6_15[15:0] = lb1d_9__out_15[15:0];
  assign out_6_16[15:0] = lb1d_9__out_16[15:0];
  assign out_6_17[15:0] = lb1d_9__out_17[15:0];
  assign out_6_18[15:0] = lb1d_9__out_18[15:0];
  assign out_6_19[15:0] = lb1d_9__out_19[15:0];

endmodule //linebuffer_U0

module Downscale (
  input  CLK,
  input [15:0] I_0_0,
  output [15:0] O,
  output  V,
  input  WE
);
  //Wire declarations for instance 'inst0' (Module linebuffer_U0)
  wire  inst0__clk;
  wire [15:0] inst0__in_0_0;
  wire [15:0] inst0__out_0_0;
  wire [15:0] inst0__out_0_1;
  wire [15:0] inst0__out_0_10;
  wire [15:0] inst0__out_0_11;
  wire [15:0] inst0__out_0_12;
  wire [15:0] inst0__out_0_13;
  wire [15:0] inst0__out_0_14;
  wire [15:0] inst0__out_0_15;
  wire [15:0] inst0__out_0_16;
  wire [15:0] inst0__out_0_17;
  wire [15:0] inst0__out_0_18;
  wire [15:0] inst0__out_0_19;
  wire [15:0] inst0__out_0_2;
  wire [15:0] inst0__out_0_3;
  wire [15:0] inst0__out_0_4;
  wire [15:0] inst0__out_0_5;
  wire [15:0] inst0__out_0_6;
  wire [15:0] inst0__out_0_7;
  wire [15:0] inst0__out_0_8;
  wire [15:0] inst0__out_0_9;
  wire [15:0] inst0__out_10_0;
  wire [15:0] inst0__out_10_1;
  wire [15:0] inst0__out_10_10;
  wire [15:0] inst0__out_10_11;
  wire [15:0] inst0__out_10_12;
  wire [15:0] inst0__out_10_13;
  wire [15:0] inst0__out_10_14;
  wire [15:0] inst0__out_10_15;
  wire [15:0] inst0__out_10_16;
  wire [15:0] inst0__out_10_17;
  wire [15:0] inst0__out_10_18;
  wire [15:0] inst0__out_10_19;
  wire [15:0] inst0__out_10_2;
  wire [15:0] inst0__out_10_3;
  wire [15:0] inst0__out_10_4;
  wire [15:0] inst0__out_10_5;
  wire [15:0] inst0__out_10_6;
  wire [15:0] inst0__out_10_7;
  wire [15:0] inst0__out_10_8;
  wire [15:0] inst0__out_10_9;
  wire [15:0] inst0__out_11_0;
  wire [15:0] inst0__out_11_1;
  wire [15:0] inst0__out_11_10;
  wire [15:0] inst0__out_11_11;
  wire [15:0] inst0__out_11_12;
  wire [15:0] inst0__out_11_13;
  wire [15:0] inst0__out_11_14;
  wire [15:0] inst0__out_11_15;
  wire [15:0] inst0__out_11_16;
  wire [15:0] inst0__out_11_17;
  wire [15:0] inst0__out_11_18;
  wire [15:0] inst0__out_11_19;
  wire [15:0] inst0__out_11_2;
  wire [15:0] inst0__out_11_3;
  wire [15:0] inst0__out_11_4;
  wire [15:0] inst0__out_11_5;
  wire [15:0] inst0__out_11_6;
  wire [15:0] inst0__out_11_7;
  wire [15:0] inst0__out_11_8;
  wire [15:0] inst0__out_11_9;
  wire [15:0] inst0__out_12_0;
  wire [15:0] inst0__out_12_1;
  wire [15:0] inst0__out_12_10;
  wire [15:0] inst0__out_12_11;
  wire [15:0] inst0__out_12_12;
  wire [15:0] inst0__out_12_13;
  wire [15:0] inst0__out_12_14;
  wire [15:0] inst0__out_12_15;
  wire [15:0] inst0__out_12_16;
  wire [15:0] inst0__out_12_17;
  wire [15:0] inst0__out_12_18;
  wire [15:0] inst0__out_12_19;
  wire [15:0] inst0__out_12_2;
  wire [15:0] inst0__out_12_3;
  wire [15:0] inst0__out_12_4;
  wire [15:0] inst0__out_12_5;
  wire [15:0] inst0__out_12_6;
  wire [15:0] inst0__out_12_7;
  wire [15:0] inst0__out_12_8;
  wire [15:0] inst0__out_12_9;
  wire [15:0] inst0__out_13_0;
  wire [15:0] inst0__out_13_1;
  wire [15:0] inst0__out_13_10;
  wire [15:0] inst0__out_13_11;
  wire [15:0] inst0__out_13_12;
  wire [15:0] inst0__out_13_13;
  wire [15:0] inst0__out_13_14;
  wire [15:0] inst0__out_13_15;
  wire [15:0] inst0__out_13_16;
  wire [15:0] inst0__out_13_17;
  wire [15:0] inst0__out_13_18;
  wire [15:0] inst0__out_13_19;
  wire [15:0] inst0__out_13_2;
  wire [15:0] inst0__out_13_3;
  wire [15:0] inst0__out_13_4;
  wire [15:0] inst0__out_13_5;
  wire [15:0] inst0__out_13_6;
  wire [15:0] inst0__out_13_7;
  wire [15:0] inst0__out_13_8;
  wire [15:0] inst0__out_13_9;
  wire [15:0] inst0__out_14_0;
  wire [15:0] inst0__out_14_1;
  wire [15:0] inst0__out_14_10;
  wire [15:0] inst0__out_14_11;
  wire [15:0] inst0__out_14_12;
  wire [15:0] inst0__out_14_13;
  wire [15:0] inst0__out_14_14;
  wire [15:0] inst0__out_14_15;
  wire [15:0] inst0__out_14_16;
  wire [15:0] inst0__out_14_17;
  wire [15:0] inst0__out_14_18;
  wire [15:0] inst0__out_14_19;
  wire [15:0] inst0__out_14_2;
  wire [15:0] inst0__out_14_3;
  wire [15:0] inst0__out_14_4;
  wire [15:0] inst0__out_14_5;
  wire [15:0] inst0__out_14_6;
  wire [15:0] inst0__out_14_7;
  wire [15:0] inst0__out_14_8;
  wire [15:0] inst0__out_14_9;
  wire [15:0] inst0__out_15_0;
  wire [15:0] inst0__out_15_1;
  wire [15:0] inst0__out_15_10;
  wire [15:0] inst0__out_15_11;
  wire [15:0] inst0__out_15_12;
  wire [15:0] inst0__out_15_13;
  wire [15:0] inst0__out_15_14;
  wire [15:0] inst0__out_15_15;
  wire [15:0] inst0__out_15_16;
  wire [15:0] inst0__out_15_17;
  wire [15:0] inst0__out_15_18;
  wire [15:0] inst0__out_15_19;
  wire [15:0] inst0__out_15_2;
  wire [15:0] inst0__out_15_3;
  wire [15:0] inst0__out_15_4;
  wire [15:0] inst0__out_15_5;
  wire [15:0] inst0__out_15_6;
  wire [15:0] inst0__out_15_7;
  wire [15:0] inst0__out_15_8;
  wire [15:0] inst0__out_15_9;
  wire [15:0] inst0__out_1_0;
  wire [15:0] inst0__out_1_1;
  wire [15:0] inst0__out_1_10;
  wire [15:0] inst0__out_1_11;
  wire [15:0] inst0__out_1_12;
  wire [15:0] inst0__out_1_13;
  wire [15:0] inst0__out_1_14;
  wire [15:0] inst0__out_1_15;
  wire [15:0] inst0__out_1_16;
  wire [15:0] inst0__out_1_17;
  wire [15:0] inst0__out_1_18;
  wire [15:0] inst0__out_1_19;
  wire [15:0] inst0__out_1_2;
  wire [15:0] inst0__out_1_3;
  wire [15:0] inst0__out_1_4;
  wire [15:0] inst0__out_1_5;
  wire [15:0] inst0__out_1_6;
  wire [15:0] inst0__out_1_7;
  wire [15:0] inst0__out_1_8;
  wire [15:0] inst0__out_1_9;
  wire [15:0] inst0__out_2_0;
  wire [15:0] inst0__out_2_1;
  wire [15:0] inst0__out_2_10;
  wire [15:0] inst0__out_2_11;
  wire [15:0] inst0__out_2_12;
  wire [15:0] inst0__out_2_13;
  wire [15:0] inst0__out_2_14;
  wire [15:0] inst0__out_2_15;
  wire [15:0] inst0__out_2_16;
  wire [15:0] inst0__out_2_17;
  wire [15:0] inst0__out_2_18;
  wire [15:0] inst0__out_2_19;
  wire [15:0] inst0__out_2_2;
  wire [15:0] inst0__out_2_3;
  wire [15:0] inst0__out_2_4;
  wire [15:0] inst0__out_2_5;
  wire [15:0] inst0__out_2_6;
  wire [15:0] inst0__out_2_7;
  wire [15:0] inst0__out_2_8;
  wire [15:0] inst0__out_2_9;
  wire [15:0] inst0__out_3_0;
  wire [15:0] inst0__out_3_1;
  wire [15:0] inst0__out_3_10;
  wire [15:0] inst0__out_3_11;
  wire [15:0] inst0__out_3_12;
  wire [15:0] inst0__out_3_13;
  wire [15:0] inst0__out_3_14;
  wire [15:0] inst0__out_3_15;
  wire [15:0] inst0__out_3_16;
  wire [15:0] inst0__out_3_17;
  wire [15:0] inst0__out_3_18;
  wire [15:0] inst0__out_3_19;
  wire [15:0] inst0__out_3_2;
  wire [15:0] inst0__out_3_3;
  wire [15:0] inst0__out_3_4;
  wire [15:0] inst0__out_3_5;
  wire [15:0] inst0__out_3_6;
  wire [15:0] inst0__out_3_7;
  wire [15:0] inst0__out_3_8;
  wire [15:0] inst0__out_3_9;
  wire [15:0] inst0__out_4_0;
  wire [15:0] inst0__out_4_1;
  wire [15:0] inst0__out_4_10;
  wire [15:0] inst0__out_4_11;
  wire [15:0] inst0__out_4_12;
  wire [15:0] inst0__out_4_13;
  wire [15:0] inst0__out_4_14;
  wire [15:0] inst0__out_4_15;
  wire [15:0] inst0__out_4_16;
  wire [15:0] inst0__out_4_17;
  wire [15:0] inst0__out_4_18;
  wire [15:0] inst0__out_4_19;
  wire [15:0] inst0__out_4_2;
  wire [15:0] inst0__out_4_3;
  wire [15:0] inst0__out_4_4;
  wire [15:0] inst0__out_4_5;
  wire [15:0] inst0__out_4_6;
  wire [15:0] inst0__out_4_7;
  wire [15:0] inst0__out_4_8;
  wire [15:0] inst0__out_4_9;
  wire [15:0] inst0__out_5_0;
  wire [15:0] inst0__out_5_1;
  wire [15:0] inst0__out_5_10;
  wire [15:0] inst0__out_5_11;
  wire [15:0] inst0__out_5_12;
  wire [15:0] inst0__out_5_13;
  wire [15:0] inst0__out_5_14;
  wire [15:0] inst0__out_5_15;
  wire [15:0] inst0__out_5_16;
  wire [15:0] inst0__out_5_17;
  wire [15:0] inst0__out_5_18;
  wire [15:0] inst0__out_5_19;
  wire [15:0] inst0__out_5_2;
  wire [15:0] inst0__out_5_3;
  wire [15:0] inst0__out_5_4;
  wire [15:0] inst0__out_5_5;
  wire [15:0] inst0__out_5_6;
  wire [15:0] inst0__out_5_7;
  wire [15:0] inst0__out_5_8;
  wire [15:0] inst0__out_5_9;
  wire [15:0] inst0__out_6_0;
  wire [15:0] inst0__out_6_1;
  wire [15:0] inst0__out_6_10;
  wire [15:0] inst0__out_6_11;
  wire [15:0] inst0__out_6_12;
  wire [15:0] inst0__out_6_13;
  wire [15:0] inst0__out_6_14;
  wire [15:0] inst0__out_6_15;
  wire [15:0] inst0__out_6_16;
  wire [15:0] inst0__out_6_17;
  wire [15:0] inst0__out_6_18;
  wire [15:0] inst0__out_6_19;
  wire [15:0] inst0__out_6_2;
  wire [15:0] inst0__out_6_3;
  wire [15:0] inst0__out_6_4;
  wire [15:0] inst0__out_6_5;
  wire [15:0] inst0__out_6_6;
  wire [15:0] inst0__out_6_7;
  wire [15:0] inst0__out_6_8;
  wire [15:0] inst0__out_6_9;
  wire [15:0] inst0__out_7_0;
  wire [15:0] inst0__out_7_1;
  wire [15:0] inst0__out_7_10;
  wire [15:0] inst0__out_7_11;
  wire [15:0] inst0__out_7_12;
  wire [15:0] inst0__out_7_13;
  wire [15:0] inst0__out_7_14;
  wire [15:0] inst0__out_7_15;
  wire [15:0] inst0__out_7_16;
  wire [15:0] inst0__out_7_17;
  wire [15:0] inst0__out_7_18;
  wire [15:0] inst0__out_7_19;
  wire [15:0] inst0__out_7_2;
  wire [15:0] inst0__out_7_3;
  wire [15:0] inst0__out_7_4;
  wire [15:0] inst0__out_7_5;
  wire [15:0] inst0__out_7_6;
  wire [15:0] inst0__out_7_7;
  wire [15:0] inst0__out_7_8;
  wire [15:0] inst0__out_7_9;
  wire [15:0] inst0__out_8_0;
  wire [15:0] inst0__out_8_1;
  wire [15:0] inst0__out_8_10;
  wire [15:0] inst0__out_8_11;
  wire [15:0] inst0__out_8_12;
  wire [15:0] inst0__out_8_13;
  wire [15:0] inst0__out_8_14;
  wire [15:0] inst0__out_8_15;
  wire [15:0] inst0__out_8_16;
  wire [15:0] inst0__out_8_17;
  wire [15:0] inst0__out_8_18;
  wire [15:0] inst0__out_8_19;
  wire [15:0] inst0__out_8_2;
  wire [15:0] inst0__out_8_3;
  wire [15:0] inst0__out_8_4;
  wire [15:0] inst0__out_8_5;
  wire [15:0] inst0__out_8_6;
  wire [15:0] inst0__out_8_7;
  wire [15:0] inst0__out_8_8;
  wire [15:0] inst0__out_8_9;
  wire [15:0] inst0__out_9_0;
  wire [15:0] inst0__out_9_1;
  wire [15:0] inst0__out_9_10;
  wire [15:0] inst0__out_9_11;
  wire [15:0] inst0__out_9_12;
  wire [15:0] inst0__out_9_13;
  wire [15:0] inst0__out_9_14;
  wire [15:0] inst0__out_9_15;
  wire [15:0] inst0__out_9_16;
  wire [15:0] inst0__out_9_17;
  wire [15:0] inst0__out_9_18;
  wire [15:0] inst0__out_9_19;
  wire [15:0] inst0__out_9_2;
  wire [15:0] inst0__out_9_3;
  wire [15:0] inst0__out_9_4;
  wire [15:0] inst0__out_9_5;
  wire [15:0] inst0__out_9_6;
  wire [15:0] inst0__out_9_7;
  wire [15:0] inst0__out_9_8;
  wire [15:0] inst0__out_9_9;
  wire  inst0__valid;
  wire  inst0__valid_chain;
  wire  inst0__wen;
  linebuffer_U0 inst0(
    .clk(inst0__clk),
    .in_0_0(inst0__in_0_0),
    .out_0_0(inst0__out_0_0),
    .out_0_1(inst0__out_0_1),
    .out_0_10(inst0__out_0_10),
    .out_0_11(inst0__out_0_11),
    .out_0_12(inst0__out_0_12),
    .out_0_13(inst0__out_0_13),
    .out_0_14(inst0__out_0_14),
    .out_0_15(inst0__out_0_15),
    .out_0_16(inst0__out_0_16),
    .out_0_17(inst0__out_0_17),
    .out_0_18(inst0__out_0_18),
    .out_0_19(inst0__out_0_19),
    .out_0_2(inst0__out_0_2),
    .out_0_3(inst0__out_0_3),
    .out_0_4(inst0__out_0_4),
    .out_0_5(inst0__out_0_5),
    .out_0_6(inst0__out_0_6),
    .out_0_7(inst0__out_0_7),
    .out_0_8(inst0__out_0_8),
    .out_0_9(inst0__out_0_9),
    .out_10_0(inst0__out_10_0),
    .out_10_1(inst0__out_10_1),
    .out_10_10(inst0__out_10_10),
    .out_10_11(inst0__out_10_11),
    .out_10_12(inst0__out_10_12),
    .out_10_13(inst0__out_10_13),
    .out_10_14(inst0__out_10_14),
    .out_10_15(inst0__out_10_15),
    .out_10_16(inst0__out_10_16),
    .out_10_17(inst0__out_10_17),
    .out_10_18(inst0__out_10_18),
    .out_10_19(inst0__out_10_19),
    .out_10_2(inst0__out_10_2),
    .out_10_3(inst0__out_10_3),
    .out_10_4(inst0__out_10_4),
    .out_10_5(inst0__out_10_5),
    .out_10_6(inst0__out_10_6),
    .out_10_7(inst0__out_10_7),
    .out_10_8(inst0__out_10_8),
    .out_10_9(inst0__out_10_9),
    .out_11_0(inst0__out_11_0),
    .out_11_1(inst0__out_11_1),
    .out_11_10(inst0__out_11_10),
    .out_11_11(inst0__out_11_11),
    .out_11_12(inst0__out_11_12),
    .out_11_13(inst0__out_11_13),
    .out_11_14(inst0__out_11_14),
    .out_11_15(inst0__out_11_15),
    .out_11_16(inst0__out_11_16),
    .out_11_17(inst0__out_11_17),
    .out_11_18(inst0__out_11_18),
    .out_11_19(inst0__out_11_19),
    .out_11_2(inst0__out_11_2),
    .out_11_3(inst0__out_11_3),
    .out_11_4(inst0__out_11_4),
    .out_11_5(inst0__out_11_5),
    .out_11_6(inst0__out_11_6),
    .out_11_7(inst0__out_11_7),
    .out_11_8(inst0__out_11_8),
    .out_11_9(inst0__out_11_9),
    .out_12_0(inst0__out_12_0),
    .out_12_1(inst0__out_12_1),
    .out_12_10(inst0__out_12_10),
    .out_12_11(inst0__out_12_11),
    .out_12_12(inst0__out_12_12),
    .out_12_13(inst0__out_12_13),
    .out_12_14(inst0__out_12_14),
    .out_12_15(inst0__out_12_15),
    .out_12_16(inst0__out_12_16),
    .out_12_17(inst0__out_12_17),
    .out_12_18(inst0__out_12_18),
    .out_12_19(inst0__out_12_19),
    .out_12_2(inst0__out_12_2),
    .out_12_3(inst0__out_12_3),
    .out_12_4(inst0__out_12_4),
    .out_12_5(inst0__out_12_5),
    .out_12_6(inst0__out_12_6),
    .out_12_7(inst0__out_12_7),
    .out_12_8(inst0__out_12_8),
    .out_12_9(inst0__out_12_9),
    .out_13_0(inst0__out_13_0),
    .out_13_1(inst0__out_13_1),
    .out_13_10(inst0__out_13_10),
    .out_13_11(inst0__out_13_11),
    .out_13_12(inst0__out_13_12),
    .out_13_13(inst0__out_13_13),
    .out_13_14(inst0__out_13_14),
    .out_13_15(inst0__out_13_15),
    .out_13_16(inst0__out_13_16),
    .out_13_17(inst0__out_13_17),
    .out_13_18(inst0__out_13_18),
    .out_13_19(inst0__out_13_19),
    .out_13_2(inst0__out_13_2),
    .out_13_3(inst0__out_13_3),
    .out_13_4(inst0__out_13_4),
    .out_13_5(inst0__out_13_5),
    .out_13_6(inst0__out_13_6),
    .out_13_7(inst0__out_13_7),
    .out_13_8(inst0__out_13_8),
    .out_13_9(inst0__out_13_9),
    .out_14_0(inst0__out_14_0),
    .out_14_1(inst0__out_14_1),
    .out_14_10(inst0__out_14_10),
    .out_14_11(inst0__out_14_11),
    .out_14_12(inst0__out_14_12),
    .out_14_13(inst0__out_14_13),
    .out_14_14(inst0__out_14_14),
    .out_14_15(inst0__out_14_15),
    .out_14_16(inst0__out_14_16),
    .out_14_17(inst0__out_14_17),
    .out_14_18(inst0__out_14_18),
    .out_14_19(inst0__out_14_19),
    .out_14_2(inst0__out_14_2),
    .out_14_3(inst0__out_14_3),
    .out_14_4(inst0__out_14_4),
    .out_14_5(inst0__out_14_5),
    .out_14_6(inst0__out_14_6),
    .out_14_7(inst0__out_14_7),
    .out_14_8(inst0__out_14_8),
    .out_14_9(inst0__out_14_9),
    .out_15_0(inst0__out_15_0),
    .out_15_1(inst0__out_15_1),
    .out_15_10(inst0__out_15_10),
    .out_15_11(inst0__out_15_11),
    .out_15_12(inst0__out_15_12),
    .out_15_13(inst0__out_15_13),
    .out_15_14(inst0__out_15_14),
    .out_15_15(inst0__out_15_15),
    .out_15_16(inst0__out_15_16),
    .out_15_17(inst0__out_15_17),
    .out_15_18(inst0__out_15_18),
    .out_15_19(inst0__out_15_19),
    .out_15_2(inst0__out_15_2),
    .out_15_3(inst0__out_15_3),
    .out_15_4(inst0__out_15_4),
    .out_15_5(inst0__out_15_5),
    .out_15_6(inst0__out_15_6),
    .out_15_7(inst0__out_15_7),
    .out_15_8(inst0__out_15_8),
    .out_15_9(inst0__out_15_9),
    .out_1_0(inst0__out_1_0),
    .out_1_1(inst0__out_1_1),
    .out_1_10(inst0__out_1_10),
    .out_1_11(inst0__out_1_11),
    .out_1_12(inst0__out_1_12),
    .out_1_13(inst0__out_1_13),
    .out_1_14(inst0__out_1_14),
    .out_1_15(inst0__out_1_15),
    .out_1_16(inst0__out_1_16),
    .out_1_17(inst0__out_1_17),
    .out_1_18(inst0__out_1_18),
    .out_1_19(inst0__out_1_19),
    .out_1_2(inst0__out_1_2),
    .out_1_3(inst0__out_1_3),
    .out_1_4(inst0__out_1_4),
    .out_1_5(inst0__out_1_5),
    .out_1_6(inst0__out_1_6),
    .out_1_7(inst0__out_1_7),
    .out_1_8(inst0__out_1_8),
    .out_1_9(inst0__out_1_9),
    .out_2_0(inst0__out_2_0),
    .out_2_1(inst0__out_2_1),
    .out_2_10(inst0__out_2_10),
    .out_2_11(inst0__out_2_11),
    .out_2_12(inst0__out_2_12),
    .out_2_13(inst0__out_2_13),
    .out_2_14(inst0__out_2_14),
    .out_2_15(inst0__out_2_15),
    .out_2_16(inst0__out_2_16),
    .out_2_17(inst0__out_2_17),
    .out_2_18(inst0__out_2_18),
    .out_2_19(inst0__out_2_19),
    .out_2_2(inst0__out_2_2),
    .out_2_3(inst0__out_2_3),
    .out_2_4(inst0__out_2_4),
    .out_2_5(inst0__out_2_5),
    .out_2_6(inst0__out_2_6),
    .out_2_7(inst0__out_2_7),
    .out_2_8(inst0__out_2_8),
    .out_2_9(inst0__out_2_9),
    .out_3_0(inst0__out_3_0),
    .out_3_1(inst0__out_3_1),
    .out_3_10(inst0__out_3_10),
    .out_3_11(inst0__out_3_11),
    .out_3_12(inst0__out_3_12),
    .out_3_13(inst0__out_3_13),
    .out_3_14(inst0__out_3_14),
    .out_3_15(inst0__out_3_15),
    .out_3_16(inst0__out_3_16),
    .out_3_17(inst0__out_3_17),
    .out_3_18(inst0__out_3_18),
    .out_3_19(inst0__out_3_19),
    .out_3_2(inst0__out_3_2),
    .out_3_3(inst0__out_3_3),
    .out_3_4(inst0__out_3_4),
    .out_3_5(inst0__out_3_5),
    .out_3_6(inst0__out_3_6),
    .out_3_7(inst0__out_3_7),
    .out_3_8(inst0__out_3_8),
    .out_3_9(inst0__out_3_9),
    .out_4_0(inst0__out_4_0),
    .out_4_1(inst0__out_4_1),
    .out_4_10(inst0__out_4_10),
    .out_4_11(inst0__out_4_11),
    .out_4_12(inst0__out_4_12),
    .out_4_13(inst0__out_4_13),
    .out_4_14(inst0__out_4_14),
    .out_4_15(inst0__out_4_15),
    .out_4_16(inst0__out_4_16),
    .out_4_17(inst0__out_4_17),
    .out_4_18(inst0__out_4_18),
    .out_4_19(inst0__out_4_19),
    .out_4_2(inst0__out_4_2),
    .out_4_3(inst0__out_4_3),
    .out_4_4(inst0__out_4_4),
    .out_4_5(inst0__out_4_5),
    .out_4_6(inst0__out_4_6),
    .out_4_7(inst0__out_4_7),
    .out_4_8(inst0__out_4_8),
    .out_4_9(inst0__out_4_9),
    .out_5_0(inst0__out_5_0),
    .out_5_1(inst0__out_5_1),
    .out_5_10(inst0__out_5_10),
    .out_5_11(inst0__out_5_11),
    .out_5_12(inst0__out_5_12),
    .out_5_13(inst0__out_5_13),
    .out_5_14(inst0__out_5_14),
    .out_5_15(inst0__out_5_15),
    .out_5_16(inst0__out_5_16),
    .out_5_17(inst0__out_5_17),
    .out_5_18(inst0__out_5_18),
    .out_5_19(inst0__out_5_19),
    .out_5_2(inst0__out_5_2),
    .out_5_3(inst0__out_5_3),
    .out_5_4(inst0__out_5_4),
    .out_5_5(inst0__out_5_5),
    .out_5_6(inst0__out_5_6),
    .out_5_7(inst0__out_5_7),
    .out_5_8(inst0__out_5_8),
    .out_5_9(inst0__out_5_9),
    .out_6_0(inst0__out_6_0),
    .out_6_1(inst0__out_6_1),
    .out_6_10(inst0__out_6_10),
    .out_6_11(inst0__out_6_11),
    .out_6_12(inst0__out_6_12),
    .out_6_13(inst0__out_6_13),
    .out_6_14(inst0__out_6_14),
    .out_6_15(inst0__out_6_15),
    .out_6_16(inst0__out_6_16),
    .out_6_17(inst0__out_6_17),
    .out_6_18(inst0__out_6_18),
    .out_6_19(inst0__out_6_19),
    .out_6_2(inst0__out_6_2),
    .out_6_3(inst0__out_6_3),
    .out_6_4(inst0__out_6_4),
    .out_6_5(inst0__out_6_5),
    .out_6_6(inst0__out_6_6),
    .out_6_7(inst0__out_6_7),
    .out_6_8(inst0__out_6_8),
    .out_6_9(inst0__out_6_9),
    .out_7_0(inst0__out_7_0),
    .out_7_1(inst0__out_7_1),
    .out_7_10(inst0__out_7_10),
    .out_7_11(inst0__out_7_11),
    .out_7_12(inst0__out_7_12),
    .out_7_13(inst0__out_7_13),
    .out_7_14(inst0__out_7_14),
    .out_7_15(inst0__out_7_15),
    .out_7_16(inst0__out_7_16),
    .out_7_17(inst0__out_7_17),
    .out_7_18(inst0__out_7_18),
    .out_7_19(inst0__out_7_19),
    .out_7_2(inst0__out_7_2),
    .out_7_3(inst0__out_7_3),
    .out_7_4(inst0__out_7_4),
    .out_7_5(inst0__out_7_5),
    .out_7_6(inst0__out_7_6),
    .out_7_7(inst0__out_7_7),
    .out_7_8(inst0__out_7_8),
    .out_7_9(inst0__out_7_9),
    .out_8_0(inst0__out_8_0),
    .out_8_1(inst0__out_8_1),
    .out_8_10(inst0__out_8_10),
    .out_8_11(inst0__out_8_11),
    .out_8_12(inst0__out_8_12),
    .out_8_13(inst0__out_8_13),
    .out_8_14(inst0__out_8_14),
    .out_8_15(inst0__out_8_15),
    .out_8_16(inst0__out_8_16),
    .out_8_17(inst0__out_8_17),
    .out_8_18(inst0__out_8_18),
    .out_8_19(inst0__out_8_19),
    .out_8_2(inst0__out_8_2),
    .out_8_3(inst0__out_8_3),
    .out_8_4(inst0__out_8_4),
    .out_8_5(inst0__out_8_5),
    .out_8_6(inst0__out_8_6),
    .out_8_7(inst0__out_8_7),
    .out_8_8(inst0__out_8_8),
    .out_8_9(inst0__out_8_9),
    .out_9_0(inst0__out_9_0),
    .out_9_1(inst0__out_9_1),
    .out_9_10(inst0__out_9_10),
    .out_9_11(inst0__out_9_11),
    .out_9_12(inst0__out_9_12),
    .out_9_13(inst0__out_9_13),
    .out_9_14(inst0__out_9_14),
    .out_9_15(inst0__out_9_15),
    .out_9_16(inst0__out_9_16),
    .out_9_17(inst0__out_9_17),
    .out_9_18(inst0__out_9_18),
    .out_9_19(inst0__out_9_19),
    .out_9_2(inst0__out_9_2),
    .out_9_3(inst0__out_9_3),
    .out_9_4(inst0__out_9_4),
    .out_9_5(inst0__out_9_5),
    .out_9_6(inst0__out_9_6),
    .out_9_7(inst0__out_9_7),
    .out_9_8(inst0__out_9_8),
    .out_9_9(inst0__out_9_9),
    .valid(inst0__valid),
    .valid_chain(inst0__valid_chain),
    .wen(inst0__wen)
  );

  //Wire declarations for instance 'inst1' (Module reduceParallel_U1)
  wire [15:0] inst1__in_data_0;
  wire [15:0] inst1__in_data_1;
  wire [15:0] inst1__in_data_10;
  wire [15:0] inst1__in_data_100;
  wire [15:0] inst1__in_data_101;
  wire [15:0] inst1__in_data_102;
  wire [15:0] inst1__in_data_103;
  wire [15:0] inst1__in_data_104;
  wire [15:0] inst1__in_data_105;
  wire [15:0] inst1__in_data_106;
  wire [15:0] inst1__in_data_107;
  wire [15:0] inst1__in_data_108;
  wire [15:0] inst1__in_data_109;
  wire [15:0] inst1__in_data_11;
  wire [15:0] inst1__in_data_110;
  wire [15:0] inst1__in_data_111;
  wire [15:0] inst1__in_data_112;
  wire [15:0] inst1__in_data_113;
  wire [15:0] inst1__in_data_114;
  wire [15:0] inst1__in_data_115;
  wire [15:0] inst1__in_data_116;
  wire [15:0] inst1__in_data_117;
  wire [15:0] inst1__in_data_118;
  wire [15:0] inst1__in_data_119;
  wire [15:0] inst1__in_data_12;
  wire [15:0] inst1__in_data_120;
  wire [15:0] inst1__in_data_121;
  wire [15:0] inst1__in_data_122;
  wire [15:0] inst1__in_data_123;
  wire [15:0] inst1__in_data_124;
  wire [15:0] inst1__in_data_125;
  wire [15:0] inst1__in_data_126;
  wire [15:0] inst1__in_data_127;
  wire [15:0] inst1__in_data_128;
  wire [15:0] inst1__in_data_129;
  wire [15:0] inst1__in_data_13;
  wire [15:0] inst1__in_data_130;
  wire [15:0] inst1__in_data_131;
  wire [15:0] inst1__in_data_132;
  wire [15:0] inst1__in_data_133;
  wire [15:0] inst1__in_data_134;
  wire [15:0] inst1__in_data_135;
  wire [15:0] inst1__in_data_136;
  wire [15:0] inst1__in_data_137;
  wire [15:0] inst1__in_data_138;
  wire [15:0] inst1__in_data_139;
  wire [15:0] inst1__in_data_14;
  wire [15:0] inst1__in_data_140;
  wire [15:0] inst1__in_data_141;
  wire [15:0] inst1__in_data_142;
  wire [15:0] inst1__in_data_143;
  wire [15:0] inst1__in_data_144;
  wire [15:0] inst1__in_data_145;
  wire [15:0] inst1__in_data_146;
  wire [15:0] inst1__in_data_147;
  wire [15:0] inst1__in_data_148;
  wire [15:0] inst1__in_data_149;
  wire [15:0] inst1__in_data_15;
  wire [15:0] inst1__in_data_150;
  wire [15:0] inst1__in_data_151;
  wire [15:0] inst1__in_data_152;
  wire [15:0] inst1__in_data_153;
  wire [15:0] inst1__in_data_154;
  wire [15:0] inst1__in_data_155;
  wire [15:0] inst1__in_data_156;
  wire [15:0] inst1__in_data_157;
  wire [15:0] inst1__in_data_158;
  wire [15:0] inst1__in_data_159;
  wire [15:0] inst1__in_data_16;
  wire [15:0] inst1__in_data_160;
  wire [15:0] inst1__in_data_161;
  wire [15:0] inst1__in_data_162;
  wire [15:0] inst1__in_data_163;
  wire [15:0] inst1__in_data_164;
  wire [15:0] inst1__in_data_165;
  wire [15:0] inst1__in_data_166;
  wire [15:0] inst1__in_data_167;
  wire [15:0] inst1__in_data_168;
  wire [15:0] inst1__in_data_169;
  wire [15:0] inst1__in_data_17;
  wire [15:0] inst1__in_data_170;
  wire [15:0] inst1__in_data_171;
  wire [15:0] inst1__in_data_172;
  wire [15:0] inst1__in_data_173;
  wire [15:0] inst1__in_data_174;
  wire [15:0] inst1__in_data_175;
  wire [15:0] inst1__in_data_176;
  wire [15:0] inst1__in_data_177;
  wire [15:0] inst1__in_data_178;
  wire [15:0] inst1__in_data_179;
  wire [15:0] inst1__in_data_18;
  wire [15:0] inst1__in_data_180;
  wire [15:0] inst1__in_data_181;
  wire [15:0] inst1__in_data_182;
  wire [15:0] inst1__in_data_183;
  wire [15:0] inst1__in_data_184;
  wire [15:0] inst1__in_data_185;
  wire [15:0] inst1__in_data_186;
  wire [15:0] inst1__in_data_187;
  wire [15:0] inst1__in_data_188;
  wire [15:0] inst1__in_data_189;
  wire [15:0] inst1__in_data_19;
  wire [15:0] inst1__in_data_190;
  wire [15:0] inst1__in_data_191;
  wire [15:0] inst1__in_data_192;
  wire [15:0] inst1__in_data_193;
  wire [15:0] inst1__in_data_194;
  wire [15:0] inst1__in_data_195;
  wire [15:0] inst1__in_data_196;
  wire [15:0] inst1__in_data_197;
  wire [15:0] inst1__in_data_198;
  wire [15:0] inst1__in_data_199;
  wire [15:0] inst1__in_data_2;
  wire [15:0] inst1__in_data_20;
  wire [15:0] inst1__in_data_200;
  wire [15:0] inst1__in_data_201;
  wire [15:0] inst1__in_data_202;
  wire [15:0] inst1__in_data_203;
  wire [15:0] inst1__in_data_204;
  wire [15:0] inst1__in_data_205;
  wire [15:0] inst1__in_data_206;
  wire [15:0] inst1__in_data_207;
  wire [15:0] inst1__in_data_208;
  wire [15:0] inst1__in_data_209;
  wire [15:0] inst1__in_data_21;
  wire [15:0] inst1__in_data_210;
  wire [15:0] inst1__in_data_211;
  wire [15:0] inst1__in_data_212;
  wire [15:0] inst1__in_data_213;
  wire [15:0] inst1__in_data_214;
  wire [15:0] inst1__in_data_215;
  wire [15:0] inst1__in_data_216;
  wire [15:0] inst1__in_data_217;
  wire [15:0] inst1__in_data_218;
  wire [15:0] inst1__in_data_219;
  wire [15:0] inst1__in_data_22;
  wire [15:0] inst1__in_data_220;
  wire [15:0] inst1__in_data_221;
  wire [15:0] inst1__in_data_222;
  wire [15:0] inst1__in_data_223;
  wire [15:0] inst1__in_data_224;
  wire [15:0] inst1__in_data_225;
  wire [15:0] inst1__in_data_226;
  wire [15:0] inst1__in_data_227;
  wire [15:0] inst1__in_data_228;
  wire [15:0] inst1__in_data_229;
  wire [15:0] inst1__in_data_23;
  wire [15:0] inst1__in_data_230;
  wire [15:0] inst1__in_data_231;
  wire [15:0] inst1__in_data_232;
  wire [15:0] inst1__in_data_233;
  wire [15:0] inst1__in_data_234;
  wire [15:0] inst1__in_data_235;
  wire [15:0] inst1__in_data_236;
  wire [15:0] inst1__in_data_237;
  wire [15:0] inst1__in_data_238;
  wire [15:0] inst1__in_data_239;
  wire [15:0] inst1__in_data_24;
  wire [15:0] inst1__in_data_240;
  wire [15:0] inst1__in_data_241;
  wire [15:0] inst1__in_data_242;
  wire [15:0] inst1__in_data_243;
  wire [15:0] inst1__in_data_244;
  wire [15:0] inst1__in_data_245;
  wire [15:0] inst1__in_data_246;
  wire [15:0] inst1__in_data_247;
  wire [15:0] inst1__in_data_248;
  wire [15:0] inst1__in_data_249;
  wire [15:0] inst1__in_data_25;
  wire [15:0] inst1__in_data_250;
  wire [15:0] inst1__in_data_251;
  wire [15:0] inst1__in_data_252;
  wire [15:0] inst1__in_data_253;
  wire [15:0] inst1__in_data_254;
  wire [15:0] inst1__in_data_255;
  wire [15:0] inst1__in_data_256;
  wire [15:0] inst1__in_data_257;
  wire [15:0] inst1__in_data_258;
  wire [15:0] inst1__in_data_259;
  wire [15:0] inst1__in_data_26;
  wire [15:0] inst1__in_data_260;
  wire [15:0] inst1__in_data_261;
  wire [15:0] inst1__in_data_262;
  wire [15:0] inst1__in_data_263;
  wire [15:0] inst1__in_data_264;
  wire [15:0] inst1__in_data_265;
  wire [15:0] inst1__in_data_266;
  wire [15:0] inst1__in_data_267;
  wire [15:0] inst1__in_data_268;
  wire [15:0] inst1__in_data_269;
  wire [15:0] inst1__in_data_27;
  wire [15:0] inst1__in_data_270;
  wire [15:0] inst1__in_data_271;
  wire [15:0] inst1__in_data_272;
  wire [15:0] inst1__in_data_273;
  wire [15:0] inst1__in_data_274;
  wire [15:0] inst1__in_data_275;
  wire [15:0] inst1__in_data_276;
  wire [15:0] inst1__in_data_277;
  wire [15:0] inst1__in_data_278;
  wire [15:0] inst1__in_data_279;
  wire [15:0] inst1__in_data_28;
  wire [15:0] inst1__in_data_280;
  wire [15:0] inst1__in_data_281;
  wire [15:0] inst1__in_data_282;
  wire [15:0] inst1__in_data_283;
  wire [15:0] inst1__in_data_284;
  wire [15:0] inst1__in_data_285;
  wire [15:0] inst1__in_data_286;
  wire [15:0] inst1__in_data_287;
  wire [15:0] inst1__in_data_288;
  wire [15:0] inst1__in_data_289;
  wire [15:0] inst1__in_data_29;
  wire [15:0] inst1__in_data_290;
  wire [15:0] inst1__in_data_291;
  wire [15:0] inst1__in_data_292;
  wire [15:0] inst1__in_data_293;
  wire [15:0] inst1__in_data_294;
  wire [15:0] inst1__in_data_295;
  wire [15:0] inst1__in_data_296;
  wire [15:0] inst1__in_data_297;
  wire [15:0] inst1__in_data_298;
  wire [15:0] inst1__in_data_299;
  wire [15:0] inst1__in_data_3;
  wire [15:0] inst1__in_data_30;
  wire [15:0] inst1__in_data_31;
  wire [15:0] inst1__in_data_32;
  wire [15:0] inst1__in_data_33;
  wire [15:0] inst1__in_data_34;
  wire [15:0] inst1__in_data_35;
  wire [15:0] inst1__in_data_36;
  wire [15:0] inst1__in_data_37;
  wire [15:0] inst1__in_data_38;
  wire [15:0] inst1__in_data_39;
  wire [15:0] inst1__in_data_4;
  wire [15:0] inst1__in_data_40;
  wire [15:0] inst1__in_data_41;
  wire [15:0] inst1__in_data_42;
  wire [15:0] inst1__in_data_43;
  wire [15:0] inst1__in_data_44;
  wire [15:0] inst1__in_data_45;
  wire [15:0] inst1__in_data_46;
  wire [15:0] inst1__in_data_47;
  wire [15:0] inst1__in_data_48;
  wire [15:0] inst1__in_data_49;
  wire [15:0] inst1__in_data_5;
  wire [15:0] inst1__in_data_50;
  wire [15:0] inst1__in_data_51;
  wire [15:0] inst1__in_data_52;
  wire [15:0] inst1__in_data_53;
  wire [15:0] inst1__in_data_54;
  wire [15:0] inst1__in_data_55;
  wire [15:0] inst1__in_data_56;
  wire [15:0] inst1__in_data_57;
  wire [15:0] inst1__in_data_58;
  wire [15:0] inst1__in_data_59;
  wire [15:0] inst1__in_data_6;
  wire [15:0] inst1__in_data_60;
  wire [15:0] inst1__in_data_61;
  wire [15:0] inst1__in_data_62;
  wire [15:0] inst1__in_data_63;
  wire [15:0] inst1__in_data_64;
  wire [15:0] inst1__in_data_65;
  wire [15:0] inst1__in_data_66;
  wire [15:0] inst1__in_data_67;
  wire [15:0] inst1__in_data_68;
  wire [15:0] inst1__in_data_69;
  wire [15:0] inst1__in_data_7;
  wire [15:0] inst1__in_data_70;
  wire [15:0] inst1__in_data_71;
  wire [15:0] inst1__in_data_72;
  wire [15:0] inst1__in_data_73;
  wire [15:0] inst1__in_data_74;
  wire [15:0] inst1__in_data_75;
  wire [15:0] inst1__in_data_76;
  wire [15:0] inst1__in_data_77;
  wire [15:0] inst1__in_data_78;
  wire [15:0] inst1__in_data_79;
  wire [15:0] inst1__in_data_8;
  wire [15:0] inst1__in_data_80;
  wire [15:0] inst1__in_data_81;
  wire [15:0] inst1__in_data_82;
  wire [15:0] inst1__in_data_83;
  wire [15:0] inst1__in_data_84;
  wire [15:0] inst1__in_data_85;
  wire [15:0] inst1__in_data_86;
  wire [15:0] inst1__in_data_87;
  wire [15:0] inst1__in_data_88;
  wire [15:0] inst1__in_data_89;
  wire [15:0] inst1__in_data_9;
  wire [15:0] inst1__in_data_90;
  wire [15:0] inst1__in_data_91;
  wire [15:0] inst1__in_data_92;
  wire [15:0] inst1__in_data_93;
  wire [15:0] inst1__in_data_94;
  wire [15:0] inst1__in_data_95;
  wire [15:0] inst1__in_data_96;
  wire [15:0] inst1__in_data_97;
  wire [15:0] inst1__in_data_98;
  wire [15:0] inst1__in_data_99;
  wire [15:0] inst1__in_identity;
  wire [15:0] inst1__out;
  reduceParallel_U1 inst1(
    .in_data_0(inst1__in_data_0),
    .in_data_1(inst1__in_data_1),
    .in_data_10(inst1__in_data_10),
    .in_data_100(inst1__in_data_100),
    .in_data_101(inst1__in_data_101),
    .in_data_102(inst1__in_data_102),
    .in_data_103(inst1__in_data_103),
    .in_data_104(inst1__in_data_104),
    .in_data_105(inst1__in_data_105),
    .in_data_106(inst1__in_data_106),
    .in_data_107(inst1__in_data_107),
    .in_data_108(inst1__in_data_108),
    .in_data_109(inst1__in_data_109),
    .in_data_11(inst1__in_data_11),
    .in_data_110(inst1__in_data_110),
    .in_data_111(inst1__in_data_111),
    .in_data_112(inst1__in_data_112),
    .in_data_113(inst1__in_data_113),
    .in_data_114(inst1__in_data_114),
    .in_data_115(inst1__in_data_115),
    .in_data_116(inst1__in_data_116),
    .in_data_117(inst1__in_data_117),
    .in_data_118(inst1__in_data_118),
    .in_data_119(inst1__in_data_119),
    .in_data_12(inst1__in_data_12),
    .in_data_120(inst1__in_data_120),
    .in_data_121(inst1__in_data_121),
    .in_data_122(inst1__in_data_122),
    .in_data_123(inst1__in_data_123),
    .in_data_124(inst1__in_data_124),
    .in_data_125(inst1__in_data_125),
    .in_data_126(inst1__in_data_126),
    .in_data_127(inst1__in_data_127),
    .in_data_128(inst1__in_data_128),
    .in_data_129(inst1__in_data_129),
    .in_data_13(inst1__in_data_13),
    .in_data_130(inst1__in_data_130),
    .in_data_131(inst1__in_data_131),
    .in_data_132(inst1__in_data_132),
    .in_data_133(inst1__in_data_133),
    .in_data_134(inst1__in_data_134),
    .in_data_135(inst1__in_data_135),
    .in_data_136(inst1__in_data_136),
    .in_data_137(inst1__in_data_137),
    .in_data_138(inst1__in_data_138),
    .in_data_139(inst1__in_data_139),
    .in_data_14(inst1__in_data_14),
    .in_data_140(inst1__in_data_140),
    .in_data_141(inst1__in_data_141),
    .in_data_142(inst1__in_data_142),
    .in_data_143(inst1__in_data_143),
    .in_data_144(inst1__in_data_144),
    .in_data_145(inst1__in_data_145),
    .in_data_146(inst1__in_data_146),
    .in_data_147(inst1__in_data_147),
    .in_data_148(inst1__in_data_148),
    .in_data_149(inst1__in_data_149),
    .in_data_15(inst1__in_data_15),
    .in_data_150(inst1__in_data_150),
    .in_data_151(inst1__in_data_151),
    .in_data_152(inst1__in_data_152),
    .in_data_153(inst1__in_data_153),
    .in_data_154(inst1__in_data_154),
    .in_data_155(inst1__in_data_155),
    .in_data_156(inst1__in_data_156),
    .in_data_157(inst1__in_data_157),
    .in_data_158(inst1__in_data_158),
    .in_data_159(inst1__in_data_159),
    .in_data_16(inst1__in_data_16),
    .in_data_160(inst1__in_data_160),
    .in_data_161(inst1__in_data_161),
    .in_data_162(inst1__in_data_162),
    .in_data_163(inst1__in_data_163),
    .in_data_164(inst1__in_data_164),
    .in_data_165(inst1__in_data_165),
    .in_data_166(inst1__in_data_166),
    .in_data_167(inst1__in_data_167),
    .in_data_168(inst1__in_data_168),
    .in_data_169(inst1__in_data_169),
    .in_data_17(inst1__in_data_17),
    .in_data_170(inst1__in_data_170),
    .in_data_171(inst1__in_data_171),
    .in_data_172(inst1__in_data_172),
    .in_data_173(inst1__in_data_173),
    .in_data_174(inst1__in_data_174),
    .in_data_175(inst1__in_data_175),
    .in_data_176(inst1__in_data_176),
    .in_data_177(inst1__in_data_177),
    .in_data_178(inst1__in_data_178),
    .in_data_179(inst1__in_data_179),
    .in_data_18(inst1__in_data_18),
    .in_data_180(inst1__in_data_180),
    .in_data_181(inst1__in_data_181),
    .in_data_182(inst1__in_data_182),
    .in_data_183(inst1__in_data_183),
    .in_data_184(inst1__in_data_184),
    .in_data_185(inst1__in_data_185),
    .in_data_186(inst1__in_data_186),
    .in_data_187(inst1__in_data_187),
    .in_data_188(inst1__in_data_188),
    .in_data_189(inst1__in_data_189),
    .in_data_19(inst1__in_data_19),
    .in_data_190(inst1__in_data_190),
    .in_data_191(inst1__in_data_191),
    .in_data_192(inst1__in_data_192),
    .in_data_193(inst1__in_data_193),
    .in_data_194(inst1__in_data_194),
    .in_data_195(inst1__in_data_195),
    .in_data_196(inst1__in_data_196),
    .in_data_197(inst1__in_data_197),
    .in_data_198(inst1__in_data_198),
    .in_data_199(inst1__in_data_199),
    .in_data_2(inst1__in_data_2),
    .in_data_20(inst1__in_data_20),
    .in_data_200(inst1__in_data_200),
    .in_data_201(inst1__in_data_201),
    .in_data_202(inst1__in_data_202),
    .in_data_203(inst1__in_data_203),
    .in_data_204(inst1__in_data_204),
    .in_data_205(inst1__in_data_205),
    .in_data_206(inst1__in_data_206),
    .in_data_207(inst1__in_data_207),
    .in_data_208(inst1__in_data_208),
    .in_data_209(inst1__in_data_209),
    .in_data_21(inst1__in_data_21),
    .in_data_210(inst1__in_data_210),
    .in_data_211(inst1__in_data_211),
    .in_data_212(inst1__in_data_212),
    .in_data_213(inst1__in_data_213),
    .in_data_214(inst1__in_data_214),
    .in_data_215(inst1__in_data_215),
    .in_data_216(inst1__in_data_216),
    .in_data_217(inst1__in_data_217),
    .in_data_218(inst1__in_data_218),
    .in_data_219(inst1__in_data_219),
    .in_data_22(inst1__in_data_22),
    .in_data_220(inst1__in_data_220),
    .in_data_221(inst1__in_data_221),
    .in_data_222(inst1__in_data_222),
    .in_data_223(inst1__in_data_223),
    .in_data_224(inst1__in_data_224),
    .in_data_225(inst1__in_data_225),
    .in_data_226(inst1__in_data_226),
    .in_data_227(inst1__in_data_227),
    .in_data_228(inst1__in_data_228),
    .in_data_229(inst1__in_data_229),
    .in_data_23(inst1__in_data_23),
    .in_data_230(inst1__in_data_230),
    .in_data_231(inst1__in_data_231),
    .in_data_232(inst1__in_data_232),
    .in_data_233(inst1__in_data_233),
    .in_data_234(inst1__in_data_234),
    .in_data_235(inst1__in_data_235),
    .in_data_236(inst1__in_data_236),
    .in_data_237(inst1__in_data_237),
    .in_data_238(inst1__in_data_238),
    .in_data_239(inst1__in_data_239),
    .in_data_24(inst1__in_data_24),
    .in_data_240(inst1__in_data_240),
    .in_data_241(inst1__in_data_241),
    .in_data_242(inst1__in_data_242),
    .in_data_243(inst1__in_data_243),
    .in_data_244(inst1__in_data_244),
    .in_data_245(inst1__in_data_245),
    .in_data_246(inst1__in_data_246),
    .in_data_247(inst1__in_data_247),
    .in_data_248(inst1__in_data_248),
    .in_data_249(inst1__in_data_249),
    .in_data_25(inst1__in_data_25),
    .in_data_250(inst1__in_data_250),
    .in_data_251(inst1__in_data_251),
    .in_data_252(inst1__in_data_252),
    .in_data_253(inst1__in_data_253),
    .in_data_254(inst1__in_data_254),
    .in_data_255(inst1__in_data_255),
    .in_data_256(inst1__in_data_256),
    .in_data_257(inst1__in_data_257),
    .in_data_258(inst1__in_data_258),
    .in_data_259(inst1__in_data_259),
    .in_data_26(inst1__in_data_26),
    .in_data_260(inst1__in_data_260),
    .in_data_261(inst1__in_data_261),
    .in_data_262(inst1__in_data_262),
    .in_data_263(inst1__in_data_263),
    .in_data_264(inst1__in_data_264),
    .in_data_265(inst1__in_data_265),
    .in_data_266(inst1__in_data_266),
    .in_data_267(inst1__in_data_267),
    .in_data_268(inst1__in_data_268),
    .in_data_269(inst1__in_data_269),
    .in_data_27(inst1__in_data_27),
    .in_data_270(inst1__in_data_270),
    .in_data_271(inst1__in_data_271),
    .in_data_272(inst1__in_data_272),
    .in_data_273(inst1__in_data_273),
    .in_data_274(inst1__in_data_274),
    .in_data_275(inst1__in_data_275),
    .in_data_276(inst1__in_data_276),
    .in_data_277(inst1__in_data_277),
    .in_data_278(inst1__in_data_278),
    .in_data_279(inst1__in_data_279),
    .in_data_28(inst1__in_data_28),
    .in_data_280(inst1__in_data_280),
    .in_data_281(inst1__in_data_281),
    .in_data_282(inst1__in_data_282),
    .in_data_283(inst1__in_data_283),
    .in_data_284(inst1__in_data_284),
    .in_data_285(inst1__in_data_285),
    .in_data_286(inst1__in_data_286),
    .in_data_287(inst1__in_data_287),
    .in_data_288(inst1__in_data_288),
    .in_data_289(inst1__in_data_289),
    .in_data_29(inst1__in_data_29),
    .in_data_290(inst1__in_data_290),
    .in_data_291(inst1__in_data_291),
    .in_data_292(inst1__in_data_292),
    .in_data_293(inst1__in_data_293),
    .in_data_294(inst1__in_data_294),
    .in_data_295(inst1__in_data_295),
    .in_data_296(inst1__in_data_296),
    .in_data_297(inst1__in_data_297),
    .in_data_298(inst1__in_data_298),
    .in_data_299(inst1__in_data_299),
    .in_data_3(inst1__in_data_3),
    .in_data_30(inst1__in_data_30),
    .in_data_31(inst1__in_data_31),
    .in_data_32(inst1__in_data_32),
    .in_data_33(inst1__in_data_33),
    .in_data_34(inst1__in_data_34),
    .in_data_35(inst1__in_data_35),
    .in_data_36(inst1__in_data_36),
    .in_data_37(inst1__in_data_37),
    .in_data_38(inst1__in_data_38),
    .in_data_39(inst1__in_data_39),
    .in_data_4(inst1__in_data_4),
    .in_data_40(inst1__in_data_40),
    .in_data_41(inst1__in_data_41),
    .in_data_42(inst1__in_data_42),
    .in_data_43(inst1__in_data_43),
    .in_data_44(inst1__in_data_44),
    .in_data_45(inst1__in_data_45),
    .in_data_46(inst1__in_data_46),
    .in_data_47(inst1__in_data_47),
    .in_data_48(inst1__in_data_48),
    .in_data_49(inst1__in_data_49),
    .in_data_5(inst1__in_data_5),
    .in_data_50(inst1__in_data_50),
    .in_data_51(inst1__in_data_51),
    .in_data_52(inst1__in_data_52),
    .in_data_53(inst1__in_data_53),
    .in_data_54(inst1__in_data_54),
    .in_data_55(inst1__in_data_55),
    .in_data_56(inst1__in_data_56),
    .in_data_57(inst1__in_data_57),
    .in_data_58(inst1__in_data_58),
    .in_data_59(inst1__in_data_59),
    .in_data_6(inst1__in_data_6),
    .in_data_60(inst1__in_data_60),
    .in_data_61(inst1__in_data_61),
    .in_data_62(inst1__in_data_62),
    .in_data_63(inst1__in_data_63),
    .in_data_64(inst1__in_data_64),
    .in_data_65(inst1__in_data_65),
    .in_data_66(inst1__in_data_66),
    .in_data_67(inst1__in_data_67),
    .in_data_68(inst1__in_data_68),
    .in_data_69(inst1__in_data_69),
    .in_data_7(inst1__in_data_7),
    .in_data_70(inst1__in_data_70),
    .in_data_71(inst1__in_data_71),
    .in_data_72(inst1__in_data_72),
    .in_data_73(inst1__in_data_73),
    .in_data_74(inst1__in_data_74),
    .in_data_75(inst1__in_data_75),
    .in_data_76(inst1__in_data_76),
    .in_data_77(inst1__in_data_77),
    .in_data_78(inst1__in_data_78),
    .in_data_79(inst1__in_data_79),
    .in_data_8(inst1__in_data_8),
    .in_data_80(inst1__in_data_80),
    .in_data_81(inst1__in_data_81),
    .in_data_82(inst1__in_data_82),
    .in_data_83(inst1__in_data_83),
    .in_data_84(inst1__in_data_84),
    .in_data_85(inst1__in_data_85),
    .in_data_86(inst1__in_data_86),
    .in_data_87(inst1__in_data_87),
    .in_data_88(inst1__in_data_88),
    .in_data_89(inst1__in_data_89),
    .in_data_9(inst1__in_data_9),
    .in_data_90(inst1__in_data_90),
    .in_data_91(inst1__in_data_91),
    .in_data_92(inst1__in_data_92),
    .in_data_93(inst1__in_data_93),
    .in_data_94(inst1__in_data_94),
    .in_data_95(inst1__in_data_95),
    .in_data_96(inst1__in_data_96),
    .in_data_97(inst1__in_data_97),
    .in_data_98(inst1__in_data_98),
    .in_data_99(inst1__in_data_99),
    .in_identity(inst1__in_identity),
    .out(inst1__out)
  );

  //Wire declarations for instance 'inst2' (Module coreir_const160)
  wire [15:0] inst2__out;
  coreir_const160 inst2(
    .out(inst2__out)
  );

  //All the connections
  assign V = inst0__valid;
  assign inst0__wen = WE;
  assign O[15:0] = inst1__out[15:0];
  assign inst1__in_identity[15:0] = inst2__out[15:0];
  assign inst0__clk = CLK;
  assign inst0__in_0_0[15:0] = I_0_0[15:0];
  assign inst1__in_data_0[15:0] = inst0__out_0_0[15:0];
  assign inst1__in_data_4[15:0] = inst0__out_0_4[15:0];
  assign inst1__in_data_5[15:0] = inst0__out_0_5[15:0];
  assign inst1__in_data_6[15:0] = inst0__out_0_6[15:0];
  assign inst1__in_data_177[15:0] = inst0__out_8_17[15:0];
  assign inst1__in_data_1[15:0] = inst0__out_0_1[15:0];
  assign inst1__in_data_2[15:0] = inst0__out_0_2[15:0];
  assign inst1__in_data_3[15:0] = inst0__out_0_3[15:0];
  assign inst1__in_data_7[15:0] = inst0__out_0_7[15:0];
  assign inst1__in_data_8[15:0] = inst0__out_0_8[15:0];
  assign inst1__in_data_9[15:0] = inst0__out_0_9[15:0];
  assign inst1__in_data_10[15:0] = inst0__out_0_10[15:0];
  assign inst1__in_data_11[15:0] = inst0__out_0_11[15:0];
  assign inst1__in_data_12[15:0] = inst0__out_0_12[15:0];
  assign inst1__in_data_13[15:0] = inst0__out_0_13[15:0];
  assign inst1__in_data_14[15:0] = inst0__out_0_14[15:0];
  assign inst1__in_data_15[15:0] = inst0__out_0_15[15:0];
  assign inst1__in_data_16[15:0] = inst0__out_0_16[15:0];
  assign inst1__in_data_17[15:0] = inst0__out_0_17[15:0];
  assign inst1__in_data_18[15:0] = inst0__out_0_18[15:0];
  assign inst1__in_data_19[15:0] = inst0__out_0_19[15:0];
  assign inst1__in_data_20[15:0] = inst0__out_1_0[15:0];
  assign inst1__in_data_21[15:0] = inst0__out_1_1[15:0];
  assign inst1__in_data_22[15:0] = inst0__out_1_2[15:0];
  assign inst1__in_data_23[15:0] = inst0__out_1_3[15:0];
  assign inst1__in_data_24[15:0] = inst0__out_1_4[15:0];
  assign inst1__in_data_25[15:0] = inst0__out_1_5[15:0];
  assign inst1__in_data_26[15:0] = inst0__out_1_6[15:0];
  assign inst1__in_data_27[15:0] = inst0__out_1_7[15:0];
  assign inst1__in_data_28[15:0] = inst0__out_1_8[15:0];
  assign inst1__in_data_29[15:0] = inst0__out_1_9[15:0];
  assign inst1__in_data_30[15:0] = inst0__out_1_10[15:0];
  assign inst1__in_data_31[15:0] = inst0__out_1_11[15:0];
  assign inst1__in_data_32[15:0] = inst0__out_1_12[15:0];
  assign inst1__in_data_33[15:0] = inst0__out_1_13[15:0];
  assign inst1__in_data_34[15:0] = inst0__out_1_14[15:0];
  assign inst1__in_data_35[15:0] = inst0__out_1_15[15:0];
  assign inst1__in_data_36[15:0] = inst0__out_1_16[15:0];
  assign inst1__in_data_37[15:0] = inst0__out_1_17[15:0];
  assign inst1__in_data_38[15:0] = inst0__out_1_18[15:0];
  assign inst1__in_data_39[15:0] = inst0__out_1_19[15:0];
  assign inst1__in_data_40[15:0] = inst0__out_2_0[15:0];
  assign inst1__in_data_41[15:0] = inst0__out_2_1[15:0];
  assign inst1__in_data_42[15:0] = inst0__out_2_2[15:0];
  assign inst1__in_data_43[15:0] = inst0__out_2_3[15:0];
  assign inst1__in_data_44[15:0] = inst0__out_2_4[15:0];
  assign inst1__in_data_45[15:0] = inst0__out_2_5[15:0];
  assign inst1__in_data_46[15:0] = inst0__out_2_6[15:0];
  assign inst1__in_data_47[15:0] = inst0__out_2_7[15:0];
  assign inst1__in_data_48[15:0] = inst0__out_2_8[15:0];
  assign inst1__in_data_49[15:0] = inst0__out_2_9[15:0];
  assign inst1__in_data_50[15:0] = inst0__out_2_10[15:0];
  assign inst1__in_data_51[15:0] = inst0__out_2_11[15:0];
  assign inst1__in_data_52[15:0] = inst0__out_2_12[15:0];
  assign inst1__in_data_53[15:0] = inst0__out_2_13[15:0];
  assign inst1__in_data_54[15:0] = inst0__out_2_14[15:0];
  assign inst1__in_data_55[15:0] = inst0__out_2_15[15:0];
  assign inst1__in_data_56[15:0] = inst0__out_2_16[15:0];
  assign inst1__in_data_57[15:0] = inst0__out_2_17[15:0];
  assign inst1__in_data_58[15:0] = inst0__out_2_18[15:0];
  assign inst1__in_data_59[15:0] = inst0__out_2_19[15:0];
  assign inst1__in_data_60[15:0] = inst0__out_3_0[15:0];
  assign inst1__in_data_61[15:0] = inst0__out_3_1[15:0];
  assign inst1__in_data_62[15:0] = inst0__out_3_2[15:0];
  assign inst1__in_data_63[15:0] = inst0__out_3_3[15:0];
  assign inst1__in_data_64[15:0] = inst0__out_3_4[15:0];
  assign inst1__in_data_65[15:0] = inst0__out_3_5[15:0];
  assign inst1__in_data_66[15:0] = inst0__out_3_6[15:0];
  assign inst1__in_data_67[15:0] = inst0__out_3_7[15:0];
  assign inst1__in_data_68[15:0] = inst0__out_3_8[15:0];
  assign inst1__in_data_69[15:0] = inst0__out_3_9[15:0];
  assign inst1__in_data_70[15:0] = inst0__out_3_10[15:0];
  assign inst1__in_data_71[15:0] = inst0__out_3_11[15:0];
  assign inst1__in_data_72[15:0] = inst0__out_3_12[15:0];
  assign inst1__in_data_73[15:0] = inst0__out_3_13[15:0];
  assign inst1__in_data_74[15:0] = inst0__out_3_14[15:0];
  assign inst1__in_data_75[15:0] = inst0__out_3_15[15:0];
  assign inst1__in_data_76[15:0] = inst0__out_3_16[15:0];
  assign inst1__in_data_77[15:0] = inst0__out_3_17[15:0];
  assign inst1__in_data_151[15:0] = inst0__out_7_11[15:0];
  assign inst1__in_data_78[15:0] = inst0__out_3_18[15:0];
  assign inst1__in_data_79[15:0] = inst0__out_3_19[15:0];
  assign inst1__in_data_80[15:0] = inst0__out_4_0[15:0];
  assign inst1__in_data_81[15:0] = inst0__out_4_1[15:0];
  assign inst1__in_data_82[15:0] = inst0__out_4_2[15:0];
  assign inst1__in_data_83[15:0] = inst0__out_4_3[15:0];
  assign inst1__in_data_84[15:0] = inst0__out_4_4[15:0];
  assign inst1__in_data_85[15:0] = inst0__out_4_5[15:0];
  assign inst1__in_data_86[15:0] = inst0__out_4_6[15:0];
  assign inst1__in_data_87[15:0] = inst0__out_4_7[15:0];
  assign inst1__in_data_88[15:0] = inst0__out_4_8[15:0];
  assign inst1__in_data_89[15:0] = inst0__out_4_9[15:0];
  assign inst1__in_data_90[15:0] = inst0__out_4_10[15:0];
  assign inst1__in_data_91[15:0] = inst0__out_4_11[15:0];
  assign inst1__in_data_92[15:0] = inst0__out_4_12[15:0];
  assign inst1__in_data_93[15:0] = inst0__out_4_13[15:0];
  assign inst1__in_data_94[15:0] = inst0__out_4_14[15:0];
  assign inst1__in_data_95[15:0] = inst0__out_4_15[15:0];
  assign inst1__in_data_96[15:0] = inst0__out_4_16[15:0];
  assign inst1__in_data_97[15:0] = inst0__out_4_17[15:0];
  assign inst1__in_data_98[15:0] = inst0__out_4_18[15:0];
  assign inst1__in_data_99[15:0] = inst0__out_4_19[15:0];
  assign inst1__in_data_100[15:0] = inst0__out_5_0[15:0];
  assign inst1__in_data_101[15:0] = inst0__out_5_1[15:0];
  assign inst1__in_data_102[15:0] = inst0__out_5_2[15:0];
  assign inst1__in_data_103[15:0] = inst0__out_5_3[15:0];
  assign inst1__in_data_104[15:0] = inst0__out_5_4[15:0];
  assign inst1__in_data_105[15:0] = inst0__out_5_5[15:0];
  assign inst1__in_data_106[15:0] = inst0__out_5_6[15:0];
  assign inst1__in_data_107[15:0] = inst0__out_5_7[15:0];
  assign inst1__in_data_108[15:0] = inst0__out_5_8[15:0];
  assign inst1__in_data_109[15:0] = inst0__out_5_9[15:0];
  assign inst1__in_data_110[15:0] = inst0__out_5_10[15:0];
  assign inst1__in_data_111[15:0] = inst0__out_5_11[15:0];
  assign inst1__in_data_112[15:0] = inst0__out_5_12[15:0];
  assign inst1__in_data_113[15:0] = inst0__out_5_13[15:0];
  assign inst1__in_data_114[15:0] = inst0__out_5_14[15:0];
  assign inst1__in_data_115[15:0] = inst0__out_5_15[15:0];
  assign inst1__in_data_116[15:0] = inst0__out_5_16[15:0];
  assign inst1__in_data_117[15:0] = inst0__out_5_17[15:0];
  assign inst1__in_data_118[15:0] = inst0__out_5_18[15:0];
  assign inst1__in_data_119[15:0] = inst0__out_5_19[15:0];
  assign inst1__in_data_120[15:0] = inst0__out_6_0[15:0];
  assign inst1__in_data_121[15:0] = inst0__out_6_1[15:0];
  assign inst1__in_data_122[15:0] = inst0__out_6_2[15:0];
  assign inst1__in_data_123[15:0] = inst0__out_6_3[15:0];
  assign inst1__in_data_124[15:0] = inst0__out_6_4[15:0];
  assign inst1__in_data_125[15:0] = inst0__out_6_5[15:0];
  assign inst1__in_data_126[15:0] = inst0__out_6_6[15:0];
  assign inst1__in_data_127[15:0] = inst0__out_6_7[15:0];
  assign inst1__in_data_128[15:0] = inst0__out_6_8[15:0];
  assign inst1__in_data_129[15:0] = inst0__out_6_9[15:0];
  assign inst1__in_data_130[15:0] = inst0__out_6_10[15:0];
  assign inst1__in_data_131[15:0] = inst0__out_6_11[15:0];
  assign inst1__in_data_132[15:0] = inst0__out_6_12[15:0];
  assign inst1__in_data_133[15:0] = inst0__out_6_13[15:0];
  assign inst1__in_data_134[15:0] = inst0__out_6_14[15:0];
  assign inst1__in_data_135[15:0] = inst0__out_6_15[15:0];
  assign inst1__in_data_136[15:0] = inst0__out_6_16[15:0];
  assign inst1__in_data_137[15:0] = inst0__out_6_17[15:0];
  assign inst1__in_data_138[15:0] = inst0__out_6_18[15:0];
  assign inst1__in_data_139[15:0] = inst0__out_6_19[15:0];
  assign inst1__in_data_140[15:0] = inst0__out_7_0[15:0];
  assign inst1__in_data_141[15:0] = inst0__out_7_1[15:0];
  assign inst1__in_data_142[15:0] = inst0__out_7_2[15:0];
  assign inst1__in_data_143[15:0] = inst0__out_7_3[15:0];
  assign inst1__in_data_144[15:0] = inst0__out_7_4[15:0];
  assign inst1__in_data_145[15:0] = inst0__out_7_5[15:0];
  assign inst1__in_data_146[15:0] = inst0__out_7_6[15:0];
  assign inst1__in_data_176[15:0] = inst0__out_8_16[15:0];
  assign inst1__in_data_147[15:0] = inst0__out_7_7[15:0];
  assign inst1__in_data_148[15:0] = inst0__out_7_8[15:0];
  assign inst1__in_data_149[15:0] = inst0__out_7_9[15:0];
  assign inst1__in_data_150[15:0] = inst0__out_7_10[15:0];
  assign inst1__in_data_154[15:0] = inst0__out_7_14[15:0];
  assign inst1__in_data_155[15:0] = inst0__out_7_15[15:0];
  assign inst1__in_data_156[15:0] = inst0__out_7_16[15:0];
  assign inst1__in_data_157[15:0] = inst0__out_7_17[15:0];
  assign inst1__in_data_158[15:0] = inst0__out_7_18[15:0];
  assign inst1__in_data_159[15:0] = inst0__out_7_19[15:0];
  assign inst1__in_data_160[15:0] = inst0__out_8_0[15:0];
  assign inst1__in_data_161[15:0] = inst0__out_8_1[15:0];
  assign inst1__in_data_162[15:0] = inst0__out_8_2[15:0];
  assign inst1__in_data_163[15:0] = inst0__out_8_3[15:0];
  assign inst1__in_data_164[15:0] = inst0__out_8_4[15:0];
  assign inst1__in_data_165[15:0] = inst0__out_8_5[15:0];
  assign inst1__in_data_166[15:0] = inst0__out_8_6[15:0];
  assign inst1__in_data_167[15:0] = inst0__out_8_7[15:0];
  assign inst1__in_data_168[15:0] = inst0__out_8_8[15:0];
  assign inst1__in_data_169[15:0] = inst0__out_8_9[15:0];
  assign inst1__in_data_170[15:0] = inst0__out_8_10[15:0];
  assign inst1__in_data_171[15:0] = inst0__out_8_11[15:0];
  assign inst1__in_data_172[15:0] = inst0__out_8_12[15:0];
  assign inst1__in_data_173[15:0] = inst0__out_8_13[15:0];
  assign inst1__in_data_174[15:0] = inst0__out_8_14[15:0];
  assign inst1__in_data_175[15:0] = inst0__out_8_15[15:0];
  assign inst1__in_data_178[15:0] = inst0__out_8_18[15:0];
  assign inst1__in_data_152[15:0] = inst0__out_7_12[15:0];
  assign inst1__in_data_153[15:0] = inst0__out_7_13[15:0];
  assign inst1__in_data_179[15:0] = inst0__out_8_19[15:0];
  assign inst1__in_data_180[15:0] = inst0__out_9_0[15:0];
  assign inst1__in_data_181[15:0] = inst0__out_9_1[15:0];
  assign inst1__in_data_182[15:0] = inst0__out_9_2[15:0];
  assign inst1__in_data_183[15:0] = inst0__out_9_3[15:0];
  assign inst1__in_data_184[15:0] = inst0__out_9_4[15:0];
  assign inst1__in_data_185[15:0] = inst0__out_9_5[15:0];
  assign inst1__in_data_186[15:0] = inst0__out_9_6[15:0];
  assign inst1__in_data_187[15:0] = inst0__out_9_7[15:0];
  assign inst1__in_data_188[15:0] = inst0__out_9_8[15:0];
  assign inst1__in_data_189[15:0] = inst0__out_9_9[15:0];
  assign inst1__in_data_190[15:0] = inst0__out_9_10[15:0];
  assign inst1__in_data_191[15:0] = inst0__out_9_11[15:0];
  assign inst1__in_data_192[15:0] = inst0__out_9_12[15:0];
  assign inst1__in_data_193[15:0] = inst0__out_9_13[15:0];
  assign inst1__in_data_194[15:0] = inst0__out_9_14[15:0];
  assign inst1__in_data_195[15:0] = inst0__out_9_15[15:0];
  assign inst1__in_data_196[15:0] = inst0__out_9_16[15:0];
  assign inst1__in_data_197[15:0] = inst0__out_9_17[15:0];
  assign inst1__in_data_198[15:0] = inst0__out_9_18[15:0];
  assign inst1__in_data_199[15:0] = inst0__out_9_19[15:0];
  assign inst1__in_data_200[15:0] = inst0__out_10_0[15:0];
  assign inst1__in_data_201[15:0] = inst0__out_10_1[15:0];
  assign inst1__in_data_202[15:0] = inst0__out_10_2[15:0];
  assign inst1__in_data_203[15:0] = inst0__out_10_3[15:0];
  assign inst1__in_data_204[15:0] = inst0__out_10_4[15:0];
  assign inst1__in_data_205[15:0] = inst0__out_10_5[15:0];
  assign inst1__in_data_206[15:0] = inst0__out_10_6[15:0];
  assign inst1__in_data_207[15:0] = inst0__out_10_7[15:0];
  assign inst1__in_data_208[15:0] = inst0__out_10_8[15:0];
  assign inst1__in_data_209[15:0] = inst0__out_10_9[15:0];
  assign inst1__in_data_210[15:0] = inst0__out_10_10[15:0];
  assign inst1__in_data_211[15:0] = inst0__out_10_11[15:0];
  assign inst1__in_data_212[15:0] = inst0__out_10_12[15:0];
  assign inst1__in_data_213[15:0] = inst0__out_10_13[15:0];
  assign inst1__in_data_214[15:0] = inst0__out_10_14[15:0];
  assign inst1__in_data_215[15:0] = inst0__out_10_15[15:0];
  assign inst1__in_data_216[15:0] = inst0__out_10_16[15:0];
  assign inst1__in_data_217[15:0] = inst0__out_10_17[15:0];
  assign inst1__in_data_218[15:0] = inst0__out_10_18[15:0];
  assign inst1__in_data_219[15:0] = inst0__out_10_19[15:0];
  assign inst1__in_data_220[15:0] = inst0__out_11_0[15:0];
  assign inst1__in_data_221[15:0] = inst0__out_11_1[15:0];
  assign inst1__in_data_222[15:0] = inst0__out_11_2[15:0];
  assign inst1__in_data_223[15:0] = inst0__out_11_3[15:0];
  assign inst1__in_data_224[15:0] = inst0__out_11_4[15:0];
  assign inst1__in_data_225[15:0] = inst0__out_11_5[15:0];
  assign inst1__in_data_226[15:0] = inst0__out_11_6[15:0];
  assign inst1__in_data_227[15:0] = inst0__out_11_7[15:0];
  assign inst1__in_data_228[15:0] = inst0__out_11_8[15:0];
  assign inst1__in_data_229[15:0] = inst0__out_11_9[15:0];
  assign inst1__in_data_230[15:0] = inst0__out_11_10[15:0];
  assign inst1__in_data_231[15:0] = inst0__out_11_11[15:0];
  assign inst1__in_data_232[15:0] = inst0__out_11_12[15:0];
  assign inst1__in_data_233[15:0] = inst0__out_11_13[15:0];
  assign inst1__in_data_234[15:0] = inst0__out_11_14[15:0];
  assign inst1__in_data_235[15:0] = inst0__out_11_15[15:0];
  assign inst1__in_data_236[15:0] = inst0__out_11_16[15:0];
  assign inst1__in_data_237[15:0] = inst0__out_11_17[15:0];
  assign inst1__in_data_238[15:0] = inst0__out_11_18[15:0];
  assign inst1__in_data_239[15:0] = inst0__out_11_19[15:0];
  assign inst1__in_data_240[15:0] = inst0__out_12_0[15:0];
  assign inst1__in_data_241[15:0] = inst0__out_12_1[15:0];
  assign inst1__in_data_242[15:0] = inst0__out_12_2[15:0];
  assign inst1__in_data_243[15:0] = inst0__out_12_3[15:0];
  assign inst1__in_data_244[15:0] = inst0__out_12_4[15:0];
  assign inst1__in_data_245[15:0] = inst0__out_12_5[15:0];
  assign inst1__in_data_246[15:0] = inst0__out_12_6[15:0];
  assign inst1__in_data_247[15:0] = inst0__out_12_7[15:0];
  assign inst1__in_data_248[15:0] = inst0__out_12_8[15:0];
  assign inst1__in_data_249[15:0] = inst0__out_12_9[15:0];
  assign inst1__in_data_250[15:0] = inst0__out_12_10[15:0];
  assign inst1__in_data_251[15:0] = inst0__out_12_11[15:0];
  assign inst1__in_data_252[15:0] = inst0__out_12_12[15:0];
  assign inst1__in_data_253[15:0] = inst0__out_12_13[15:0];
  assign inst1__in_data_254[15:0] = inst0__out_12_14[15:0];
  assign inst1__in_data_255[15:0] = inst0__out_12_15[15:0];
  assign inst1__in_data_256[15:0] = inst0__out_12_16[15:0];
  assign inst1__in_data_257[15:0] = inst0__out_12_17[15:0];
  assign inst1__in_data_258[15:0] = inst0__out_12_18[15:0];
  assign inst1__in_data_259[15:0] = inst0__out_12_19[15:0];
  assign inst1__in_data_260[15:0] = inst0__out_13_0[15:0];
  assign inst1__in_data_261[15:0] = inst0__out_13_1[15:0];
  assign inst1__in_data_262[15:0] = inst0__out_13_2[15:0];
  assign inst1__in_data_263[15:0] = inst0__out_13_3[15:0];
  assign inst1__in_data_264[15:0] = inst0__out_13_4[15:0];
  assign inst1__in_data_265[15:0] = inst0__out_13_5[15:0];
  assign inst1__in_data_266[15:0] = inst0__out_13_6[15:0];
  assign inst1__in_data_267[15:0] = inst0__out_13_7[15:0];
  assign inst1__in_data_268[15:0] = inst0__out_13_8[15:0];
  assign inst1__in_data_269[15:0] = inst0__out_13_9[15:0];
  assign inst1__in_data_270[15:0] = inst0__out_13_10[15:0];
  assign inst1__in_data_271[15:0] = inst0__out_13_11[15:0];
  assign inst1__in_data_272[15:0] = inst0__out_13_12[15:0];
  assign inst1__in_data_273[15:0] = inst0__out_13_13[15:0];
  assign inst1__in_data_274[15:0] = inst0__out_13_14[15:0];
  assign inst1__in_data_275[15:0] = inst0__out_13_15[15:0];
  assign inst1__in_data_276[15:0] = inst0__out_13_16[15:0];
  assign inst1__in_data_277[15:0] = inst0__out_13_17[15:0];
  assign inst1__in_data_278[15:0] = inst0__out_13_18[15:0];
  assign inst1__in_data_279[15:0] = inst0__out_13_19[15:0];
  assign inst1__in_data_280[15:0] = inst0__out_14_0[15:0];
  assign inst1__in_data_281[15:0] = inst0__out_14_1[15:0];
  assign inst1__in_data_282[15:0] = inst0__out_14_2[15:0];
  assign inst1__in_data_283[15:0] = inst0__out_14_3[15:0];
  assign inst1__in_data_284[15:0] = inst0__out_14_4[15:0];
  assign inst1__in_data_285[15:0] = inst0__out_14_5[15:0];
  assign inst1__in_data_286[15:0] = inst0__out_14_6[15:0];
  assign inst1__in_data_287[15:0] = inst0__out_14_7[15:0];
  assign inst1__in_data_288[15:0] = inst0__out_14_8[15:0];
  assign inst1__in_data_289[15:0] = inst0__out_14_9[15:0];
  assign inst1__in_data_290[15:0] = inst0__out_14_10[15:0];
  assign inst1__in_data_291[15:0] = inst0__out_14_11[15:0];
  assign inst1__in_data_292[15:0] = inst0__out_14_12[15:0];
  assign inst1__in_data_293[15:0] = inst0__out_14_13[15:0];
  assign inst1__in_data_294[15:0] = inst0__out_14_14[15:0];
  assign inst1__in_data_295[15:0] = inst0__out_14_15[15:0];
  assign inst1__in_data_296[15:0] = inst0__out_14_16[15:0];
  assign inst1__in_data_297[15:0] = inst0__out_14_17[15:0];
  assign inst1__in_data_298[15:0] = inst0__out_14_18[15:0];
  assign inst1__in_data_299[15:0] = inst0__out_14_19[15:0];

endmodule //Downscale
